module top( clk_1 , clk_2 , clk_3 , clk_4 , clk_5 , clk_6 , clk_7 , clk_8 , N1 , N101 , N106 , N111 , N116 , N121 , N126 , N13 , N130 , N135 , N138 , N143 , N146 , N149 , N152 , N153 , N156 , N159 , N165 , N17 , N171 , N177 , N183 , N189 , N195 , N201 , N207 , N210 , N219 , N228 , N237 , N246 , N255 , N259 , N26 , N260 , N261 , N267 , N268 , N29 , N36 , N42 , N51 , N55 , N59 , N68 , N72 , N73 , N74 , N75 , N8 , N80 , N85 , N86 , N87 , N88 , N89 , N90 , N91 , N96 , N388 , N389 , N390 , N391 , N418 , N419 , N420 , N421 , N422 , N423 , N446 , N447 , N448 , N449 , N450 , N767 , N768 , N850 , N863 , N864 , N865 , N866 , N874 , N878 , N879 , N880 );

input N1 , N101 , N106 , N111 , N116 , N121 , N126 , N13 , N130 , N135 , N138 , N143 , N146 , N149 , N152 , N153 , N156 , N159 , N165 , N17 , N171 , N177 , N183 , N189 , N195 , N201 , N207 , N210 , N219 , N228 , N237 , N246 , N255 , N259 , N26 , N260 , N261 , N267 , N268 , N29 , N36 , N42 , N51 , N55 , N59 , N68 , N72 , N73 , N74 , N75 , N8 , N80 , N85 , N86 , N87 , N88 , N89 , N90 , N91 , N96 ;
output N388 , N389 , N390 , N391 , N418 , N419 , N420 , N421 , N422 , N423 , N446 , N447 , N448 , N449 , N450 , N767 , N768 , N850 , N863 , N864 , N865 , N866 , N874 , N878 , N879 , N880 ;
wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , buf_N101_splitterN101ton102n316_1 , buf_N111_splitterN111ton105n207_1 , buf_N116_splitterN116ton105n190_1 , buf_N126_splitterN126ton100n163_2 , buf_N126_splitterN126ton100n163_1 , buf_N130_splitterN130ton90n121_1 , buf_N138_splitterN138ton291n283_2 , buf_N138_splitterN138ton291n283_1 , buf_N143_splitterfromN143_4 , buf_N143_splitterfromN143_3 , buf_N143_splitterfromN143_2 , buf_N143_splitterfromN143_1 , buf_N146_splitterfromN146_3 , buf_N146_splitterfromN146_2 , buf_N146_splitterfromN146_1 , buf_N149_splitterfromN149_4 , buf_N149_splitterfromN149_3 , buf_N149_splitterfromN149_2 , buf_N149_splitterfromN149_1 , buf_N152_n291_3 , buf_N152_n291_2 , buf_N152_n291_1 , buf_N153_splitterfromN153_4 , buf_N153_splitterfromN153_3 , buf_N153_splitterfromN153_2 , buf_N153_splitterfromN153_1 , buf_N207_splitterfromN207_1 , buf_N219_splitterN219ton171n325_8 , buf_N219_splitterN219ton171n325_7 , buf_N219_splitterN219ton171n325_6 , buf_N219_splitterN219ton171n325_5 , buf_N219_splitterN219ton171n325_4 , buf_N219_splitterN219ton171n325_3 , buf_N219_splitterN219ton171n325_2 , buf_N219_splitterN219ton171n325_1 , buf_N228_splitterN228ton173n342_7 , buf_N228_splitterN228ton173n342_6 , buf_N228_splitterN228ton173n342_5 , buf_N228_splitterN228ton173n342_4 , buf_N228_splitterN228ton173n342_3 , buf_N228_splitterN228ton173n342_2 , buf_N228_splitterN228ton173n342_1 , buf_N237_splitterN237ton174n328_6 , buf_N237_splitterN237ton174n328_5 , buf_N237_splitterN237ton174n328_4 , buf_N237_splitterN237ton174n328_3 , buf_N237_splitterN237ton174n328_2 , buf_N237_splitterN237ton174n328_1 , buf_N246_splitterN246ton175n359_5 , buf_N246_splitterN246ton175n359_4 , buf_N246_splitterN246ton175n359_3 , buf_N246_splitterN246ton175n359_2 , buf_N246_splitterN246ton175n359_1 , buf_N260_n254_1 , buf_N261_splitterN261ton201n170_6 , buf_N261_splitterN261ton201n170_5 , buf_N261_splitterN261ton201n170_4 , buf_N261_splitterN261ton201n170_3 , buf_N261_splitterN261ton201n170_2 , buf_N261_splitterN261ton201n170_1 , buf_N268_splitterN268ton265n331_1 , buf_N55_splitterN55ton82n263_1 , buf_N73_n177_1 , buf_N74_n87_2 , buf_N74_n87_1 , buf_N80_splitterN80ton149n76_1 , buf_N89_n89_1 , buf_N90_n79_1 , buf_N91_splitterN91ton93n345_4 , buf_N91_splitterN91ton93n345_3 , buf_N91_splitterN91ton93n345_2 , buf_N91_splitterN91ton93n345_1 , buf_N96_splitterN96ton90n360_2 , buf_N96_splitterN96ton90n360_1 , buf_n62_N388_16 , buf_n62_N388_15 , buf_n62_N388_14 , buf_n62_N388_13 , buf_n62_N388_12 , buf_n62_N388_11 , buf_n62_N388_10 , buf_n62_N388_9 , buf_n62_N388_8 , buf_n62_N388_7 , buf_n62_N388_6 , buf_n62_N388_5 , buf_n62_N388_4 , buf_n62_N388_3 , buf_n62_N388_2 , buf_n62_N388_1 , buf_n63_splitterfromn63_1 , buf_n64_N389_15 , buf_n64_N389_14 , buf_n64_N389_13 , buf_n64_N389_12 , buf_n64_N389_11 , buf_n64_N389_10 , buf_n64_N389_9 , buf_n64_N389_8 , buf_n64_N389_7 , buf_n64_N389_6 , buf_n64_N389_5 , buf_n64_N389_4 , buf_n64_N389_3 , buf_n64_N389_2 , buf_n64_N389_1 , buf_n65_splittern65ton72N390_13 , buf_n65_splittern65ton72N390_12 , buf_n65_splittern65ton72N390_11 , buf_n65_splittern65ton72N390_10 , buf_n65_splittern65ton72N390_9 , buf_n65_splittern65ton72N390_8 , buf_n65_splittern65ton72N390_7 , buf_n65_splittern65ton72N390_6 , buf_n65_splittern65ton72N390_5 , buf_n65_splittern65ton72N390_4 , buf_n65_splittern65ton72N390_3 , buf_n65_splittern65ton72N390_2 , buf_n65_splittern65ton72N390_1 , buf_n66_N391_19 , buf_n66_N391_18 , buf_n66_N391_17 , buf_n66_N391_16 , buf_n66_N391_15 , buf_n66_N391_14 , buf_n66_N391_13 , buf_n66_N391_12 , buf_n66_N391_11 , buf_n66_N391_10 , buf_n66_N391_9 , buf_n66_N391_8 , buf_n66_N391_7 , buf_n66_N391_6 , buf_n66_N391_5 , buf_n66_N391_4 , buf_n66_N391_3 , buf_n66_N391_2 , buf_n66_N391_1 , buf_n69_N418_16 , buf_n69_N418_15 , buf_n69_N418_14 , buf_n69_N418_13 , buf_n69_N418_12 , buf_n69_N418_11 , buf_n69_N418_10 , buf_n69_N418_9 , buf_n69_N418_8 , buf_n69_N418_7 , buf_n69_N418_6 , buf_n69_N418_5 , buf_n69_N418_4 , buf_n69_N418_3 , buf_n69_N418_2 , buf_n69_N418_1 , buf_n71_splitterfromn71_14 , buf_n71_splitterfromn71_13 , buf_n71_splitterfromn71_12 , buf_n71_splitterfromn71_11 , buf_n71_splitterfromn71_10 , buf_n71_splitterfromn71_9 , buf_n71_splitterfromn71_8 , buf_n71_splitterfromn71_7 , buf_n71_splitterfromn71_6 , buf_n71_splitterfromn71_5 , buf_n71_splitterfromn71_4 , buf_n71_splitterfromn71_3 , buf_n71_splitterfromn71_2 , buf_n71_splitterfromn71_1 , buf_n74_N420_15 , buf_n74_N420_14 , buf_n74_N420_13 , buf_n74_N420_12 , buf_n74_N420_11 , buf_n74_N420_10 , buf_n74_N420_9 , buf_n74_N420_8 , buf_n74_N420_7 , buf_n74_N420_6 , buf_n74_N420_5 , buf_n74_N420_4 , buf_n74_N420_3 , buf_n74_N420_2 , buf_n74_N420_1 , buf_n75_splitterfromn75_1 , buf_n76_N421_15 , buf_n76_N421_14 , buf_n76_N421_13 , buf_n76_N421_12 , buf_n76_N421_11 , buf_n76_N421_10 , buf_n76_N421_9 , buf_n76_N421_8 , buf_n76_N421_7 , buf_n76_N421_6 , buf_n76_N421_5 , buf_n76_N421_4 , buf_n76_N421_3 , buf_n76_N421_2 , buf_n76_N421_1 , buf_n77_N422_15 , buf_n77_N422_14 , buf_n77_N422_13 , buf_n77_N422_12 , buf_n77_N422_11 , buf_n77_N422_10 , buf_n77_N422_9 , buf_n77_N422_8 , buf_n77_N422_7 , buf_n77_N422_6 , buf_n77_N422_5 , buf_n77_N422_4 , buf_n77_N422_3 , buf_n77_N422_2 , buf_n77_N422_1 , buf_n79_N423_18 , buf_n79_N423_17 , buf_n79_N423_16 , buf_n79_N423_15 , buf_n79_N423_14 , buf_n79_N423_13 , buf_n79_N423_12 , buf_n79_N423_11 , buf_n79_N423_10 , buf_n79_N423_9 , buf_n79_N423_8 , buf_n79_N423_7 , buf_n79_N423_6 , buf_n79_N423_5 , buf_n79_N423_4 , buf_n79_N423_3 , buf_n79_N423_2 , buf_n79_N423_1 , buf_n84_n85_1 , buf_n85_N448_16 , buf_n85_N448_15 , buf_n85_N448_14 , buf_n85_N448_13 , buf_n85_N448_12 , buf_n85_N448_11 , buf_n85_N448_10 , buf_n85_N448_9 , buf_n85_N448_8 , buf_n85_N448_7 , buf_n85_N448_6 , buf_n85_N448_5 , buf_n85_N448_4 , buf_n85_N448_3 , buf_n85_N448_2 , buf_n85_N448_1 , buf_n88_N449_16 , buf_n88_N449_15 , buf_n88_N449_14 , buf_n88_N449_13 , buf_n88_N449_12 , buf_n88_N449_11 , buf_n88_N449_10 , buf_n88_N449_9 , buf_n88_N449_8 , buf_n88_N449_7 , buf_n88_N449_6 , buf_n88_N449_5 , buf_n88_N449_4 , buf_n88_N449_3 , buf_n88_N449_2 , buf_n88_N449_1 , buf_n89_N450_18 , buf_n89_N450_17 , buf_n89_N450_16 , buf_n89_N450_15 , buf_n89_N450_14 , buf_n89_N450_13 , buf_n89_N450_12 , buf_n89_N450_11 , buf_n89_N450_10 , buf_n89_N450_9 , buf_n89_N450_8 , buf_n89_N450_7 , buf_n89_N450_6 , buf_n89_N450_5 , buf_n89_N450_4 , buf_n89_N450_3 , buf_n89_N450_2 , buf_n89_N450_1 , buf_n116_N767_10 , buf_n116_N767_9 , buf_n116_N767_8 , buf_n116_N767_7 , buf_n116_N767_6 , buf_n116_N767_5 , buf_n116_N767_4 , buf_n116_N767_3 , buf_n116_N767_2 , buf_n116_N767_1 , buf_n143_N768_12 , buf_n143_N768_11 , buf_n143_N768_10 , buf_n143_N768_9 , buf_n143_N768_8 , buf_n143_N768_7 , buf_n143_N768_6 , buf_n143_N768_5 , buf_n143_N768_4 , buf_n143_N768_3 , buf_n143_N768_2 , buf_n143_N768_1 , buf_n181_n183_1 , buf_n183_n184_2 , buf_n183_n184_1 , buf_n184_n185_2 , buf_n184_n185_1 , buf_n188_N850_9 , buf_n188_N850_8 , buf_n188_N850_7 , buf_n188_N850_6 , buf_n188_N850_5 , buf_n188_N850_4 , buf_n188_N850_3 , buf_n188_N850_2 , buf_n188_N850_1 , buf_n224_n225_2 , buf_n224_n225_1 , buf_n226_n227_1 , buf_n227_N863_5 , buf_n227_N863_4 , buf_n227_N863_3 , buf_n227_N863_2 , buf_n227_N863_1 , buf_n238_n239_1 , buf_n239_n240_2 , buf_n239_n240_1 , buf_n240_n241_2 , buf_n240_n241_1 , buf_n241_n242_2 , buf_n241_n242_1 , buf_n243_n244_1 , buf_n244_N864_6 , buf_n244_N864_5 , buf_n244_N864_4 , buf_n244_N864_3 , buf_n244_N864_2 , buf_n244_N864_1 , buf_n256_n257_2 , buf_n256_n257_1 , buf_n257_n258_2 , buf_n257_n258_1 , buf_n258_n259_1 , buf_n260_n261_1 , buf_n261_N865_8 , buf_n261_N865_7 , buf_n261_N865_6 , buf_n261_N865_5 , buf_n261_N865_4 , buf_n261_N865_3 , buf_n261_N865_2 , buf_n261_N865_1 , buf_n271_splittern271ton328n306_3 , buf_n271_splittern271ton328n306_2 , buf_n271_splittern271ton328n306_1 , buf_n272_splitterfromn272_3 , buf_n272_splitterfromn272_2 , buf_n272_splitterfromn272_1 , buf_n279_splittern279ton343n304_2 , buf_n279_splittern279ton343n304_1 , buf_n280_splitterfromn280_3 , buf_n280_splitterfromn280_2 , buf_n280_splitterfromn280_1 , buf_n287_splittern287ton358n302_1 , buf_n288_splitterfromn288_2 , buf_n288_splitterfromn288_1 , buf_n291_n292_1 , buf_n295_splittern295ton313n300_1 , buf_n296_splitterfromn296_1 , buf_n306_N866_1 , buf_n317_n318_1 , buf_n318_n319_4 , buf_n318_n319_3 , buf_n318_n319_2 , buf_n318_n319_1 , buf_n319_n320_1 , buf_n321_N874_4 , buf_n321_N874_3 , buf_n321_N874_2 , buf_n321_N874_1 , buf_n332_n333_1 , buf_n333_n334_5 , buf_n333_n334_4 , buf_n333_n334_3 , buf_n333_n334_2 , buf_n333_n334_1 , buf_n334_n335_1 , buf_n335_n336_2 , buf_n335_n336_1 , buf_n348_n349_5 , buf_n348_n349_4 , buf_n348_n349_3 , buf_n348_n349_2 , buf_n348_n349_1 , buf_n349_n350_2 , buf_n349_n350_1 , buf_n350_n351_1 , buf_n351_N879_1 , buf_n362_n363_1 , buf_n363_n364_4 , buf_n363_n364_3 , buf_n363_n364_2 , buf_n363_n364_1 , buf_n364_n365_1 , buf_n365_n366_1 , buf_n366_N880_3 , buf_n366_N880_2 , buf_n366_N880_1 , buf_splitterN1ton70n147_n147_3 , buf_splitterN1ton70n147_n147_2 , buf_splitterN1ton70n147_n147_1 , buf_splitterN101ton102n316_splitterN101ton281n316_3 , buf_splitterN101ton102n316_splitterN101ton281n316_2 , buf_splitterN101ton102n316_splitterN101ton281n316_1 , buf_splitterN106ton102n222_splitterN106ton289n222_3 , buf_splitterN106ton102n222_splitterN106ton289n222_2 , buf_splitterN106ton102n222_splitterN106ton289n222_1 , buf_splitterN106ton289n222_n222_1 , buf_splitterN111ton105n207_n207_3 , buf_splitterN111ton105n207_n207_2 , buf_splitterN111ton105n207_n207_1 , buf_splitterN116ton105n190_n190_3 , buf_splitterN116ton105n190_n190_2 , buf_splitterN116ton105n190_n190_1 , buf_splitterN121ton182n196_n196_3 , buf_splitterN121ton182n196_n196_2 , buf_splitterN121ton182n196_n196_1 , buf_splitterN126ton100n163_n163_1 , buf_splitterfromN13_n68_1 , buf_splitterfromN146_n189_1 , buf_splitterN159ton117n272_splitterN159ton330n272_4 , buf_splitterN159ton117n272_splitterN159ton330n272_3 , buf_splitterN159ton117n272_splitterN159ton330n272_2 , buf_splitterN159ton117n272_splitterN159ton330n272_1 , buf_splitterN159ton330n272_splitterN159ton271n272_3 , buf_splitterN159ton330n272_splitterN159ton271n272_2 , buf_splitterN159ton330n272_splitterN159ton271n272_1 , buf_splitterN165ton129n280_splitterN165ton346n280_5 , buf_splitterN165ton129n280_splitterN165ton346n280_4 , buf_splitterN165ton129n280_splitterN165ton346n280_3 , buf_splitterN165ton129n280_splitterN165ton346n280_2 , buf_splitterN165ton129n280_splitterN165ton346n280_1 , buf_splitterN165ton346n280_splitterN165ton279n280_2 , buf_splitterN165ton346n280_splitterN165ton279n280_1 , buf_splitterN171ton132n288_splitterN171ton361n288_4 , buf_splitterN171ton132n288_splitterN171ton361n288_3 , buf_splitterN171ton132n288_splitterN171ton361n288_2 , buf_splitterN171ton132n288_splitterN171ton361n288_1 , buf_splitterN171ton361n288_splitterN171ton287n288_2 , buf_splitterN171ton361n288_splitterN171ton287n288_1 , buf_splitterN177ton117n296_splitterN177ton315n296_3 , buf_splitterN177ton117n296_splitterN177ton315n296_2 , buf_splitterN177ton117n296_splitterN177ton315n296_1 , buf_splitterN177ton315n296_splitterN177ton295n296_3 , buf_splitterN177ton315n296_splitterN177ton295n296_2 , buf_splitterN177ton315n296_splitterN177ton295n296_1 , buf_splitterN183ton132n212_splitterN183ton221n212_4 , buf_splitterN183ton132n212_splitterN183ton221n212_3 , buf_splitterN183ton132n212_splitterN183ton221n212_2 , buf_splitterN183ton132n212_splitterN183ton221n212_1 , buf_splitterN183ton221n212_splitterN183ton211n212_2 , buf_splitterN183ton221n212_splitterN183ton211n212_1 , buf_splitterN189ton123n194_splitterN189ton236n194_2 , buf_splitterN189ton123n194_splitterN189ton236n194_1 , buf_splitterN189ton236n194_splitterN189ton193n194_3 , buf_splitterN189ton236n194_splitterN189ton193n194_2 , buf_splitterN189ton236n194_splitterN189ton193n194_1 , buf_splitterN195ton123n200_splitterN195ton253n200_2 , buf_splitterN195ton123n200_splitterN195ton253n200_1 , buf_splitterN195ton253n200_splitterN195ton199n200_2 , buf_splitterN195ton253n200_splitterN195ton199n200_1 , buf_splitterN201ton129n167_splitterN201ton180n167_2 , buf_splitterN201ton129n167_splitterN201ton180n167_1 , buf_splitterN201ton180n167_splitterN201ton166n167_2 , buf_splitterN201ton180n167_splitterN201ton166n167_1 , buf_splitterN210ton182n345_splitterN210ton316n345_3 , buf_splitterN210ton182n345_splitterN210ton316n345_2 , buf_splitterN210ton182n345_splitterN210ton316n345_1 , buf_splitterN219ton171n325_splitterN219ton249n325_1 , buf_splitterN219ton249n325_splitterN219ton232n325_1 , buf_splitterN219ton232n325_splitterN219ton217n325_1 , buf_splitterN219ton217n325_splitterN219ton355n325_1 , buf_splitterN219ton355n325_splitterN219ton340n325_1 , buf_splitterN219ton340n325_n325_2 , buf_splitterN219ton340n325_n325_1 , buf_splitterN228ton250n342_splitterN228ton233n342_1 , buf_splitterN228ton218n342_splitterN228ton309n342_1 , buf_splitterN237ton174n328_splitterN237ton251n328_1 , buf_splitterN268ton265n331_splitterN268ton152n331_1 , buf_splitterN268ton152n331_n331_2 , buf_splitterN268ton152n331_n331_1 , buf_splitterN51ton81n275_n275_2 , buf_splitterN51ton81n275_n275_1 , buf_splitterN55ton82n263_splitterN55ton151n263_1 , buf_splitterfromN8_n267_2 , buf_splitterfromN8_n267_1 , buf_splitterN80ton149n76_splitterN80ton64n76_1 , buf_splitterN96ton90n360_splitterN96ton273n360_2 , buf_splitterN96ton90n360_splitterN96ton273n360_1 , buf_splitterN96ton273n360_n360_1 , buf_splitterfromn61_n62_1 , buf_splittern65ton72N390_N390_1 , buf_splittern67ton160n69_n69_1 , buf_splitterfromn70_n71_1 , buf_splitterfromn73_n74_1 , buf_splittern81ton145N447_N447_17 , buf_splittern81ton145N447_N447_16 , buf_splittern81ton145N447_N447_15 , buf_splittern81ton145N447_N447_14 , buf_splittern81ton145N447_N447_13 , buf_splittern81ton145N447_N447_12 , buf_splittern81ton145N447_N447_11 , buf_splittern81ton145N447_N447_10 , buf_splittern81ton145N447_N447_9 , buf_splittern81ton145N447_N447_8 , buf_splittern81ton145N447_N447_7 , buf_splittern81ton145N447_N447_6 , buf_splittern81ton145N447_N447_5 , buf_splittern81ton145N447_N447_4 , buf_splittern81ton145N447_N447_3 , buf_splittern81ton145N447_N447_2 , buf_splittern81ton145N447_N447_1 , buf_splittern152ton164n210_n210_1 , buf_splittern193ton228n206_n206_1 , buf_splittern199ton245n204_n204_1 , buf_splittern211ton213n298_n298_2 , buf_splittern211ton213n298_n298_1 , buf_splitterfromn212_n297_1 , buf_splittern271ton328n306_n306_4 , buf_splittern271ton328n306_n306_3 , buf_splittern271ton328n306_n306_2 , buf_splittern271ton328n306_n306_1 , buf_splitterfromn272_n305_4 , buf_splitterfromn272_n305_3 , buf_splitterfromn272_n305_2 , buf_splitterfromn272_n305_1 , buf_splittern279ton337n304_n304_3 , buf_splittern279ton337n304_n304_2 , buf_splittern279ton337n304_n304_1 , buf_splitterfromn280_n303_2 , buf_splitterfromn280_n303_1 , buf_splittern287ton352n302_n302_2 , buf_splittern287ton352n302_n302_1 , buf_splitterfromn288_n301_2 , buf_splitterfromn288_n301_1 , buf_splittern295ton313n300_n300_2 , buf_splittern295ton313n300_n300_1 , buf_splitterfromn296_n299_2 , buf_splitterfromn296_n299_1 , buf_splitterfromn307_n310_1 , buf_splittern322ton327n324_splittern322ton323n324_1 , splitterN1ton70n147 , splitterN101ton102n316 , splitterN101ton281n316 , splitterN106ton102n222 , splitterN106ton289n222 , splitterN111ton105n207 , splitterN116ton105n190 , splitterN121ton182n196 , splitterN126ton100n163 , splitterfromN13 , splitterN130ton90n121 , splitterN130ton120n121 , splitterfromN135 , splitterN138ton291n283 , splitterfromN143 , splitterfromN146 , splitterfromN149 , splitterfromN153 , splitterN159ton117n272 , splitterN159ton330n272 , splitterN159ton271n272 , splitterN165ton129n280 , splitterN165ton346n280 , splitterN165ton279n280 , splitterN17ton153n283 , splitterN17ton68n283 , splitterN17ton146n283 , splitterN171ton132n288 , splitterN171ton361n288 , splitterN171ton287n288 , splitterN177ton117n296 , splitterN177ton315n296 , splitterN177ton295n296 , splitterN183ton132n212 , splitterN183ton221n212 , splitterN183ton211n212 , splitterN189ton123n194 , splitterN189ton236n194 , splitterN189ton193n194 , splitterN195ton123n200 , splitterN195ton253n200 , splitterN195ton199n200 , splitterN201ton129n167 , splitterN201ton180n167 , splitterN201ton166n167 , splitterfromN207 , splitterN210ton182n345 , splitterN210ton316n345 , splitterN210ton222n345 , splitterN219ton171n325 , splitterN219ton249n325 , splitterN219ton232n325 , splitterN219ton217n325 , splitterN219ton355n325 , splitterN219ton340n325 , splitterN228ton173n342 , splitterN228ton250n342 , splitterN228ton233n342 , splitterN228ton218n342 , splitterN228ton309n342 , splitterN228ton357n342 , splitterN228ton327n342 , splitterN237ton174n328 , splitterN237ton251n328 , splitterN237ton234n328 , splitterN237ton219n328 , splitterN237ton313n328 , splitterN237ton358n328 , splitterN237ton343n328 , splitterN246ton175n359 , splitterN246ton235n359 , splitterN246ton314n359 , splitterN255ton181n254 , splitterN261ton201n170 , splitterN261ton169n170 , splitterN268ton265n331 , splitterN268ton152n331 , splitterN29ton61n84 , splitterfromN36 , splitterN42ton176n77 , splitterN42ton153n77 , splitterN42ton158n77 , splitterN42ton62n77 , splitterN51ton159n275 , splitterN51ton81n275 , splitterN55ton82n263 , splitterN55ton151n263 , splitterN59ton144n75 , splitterN59ton73n75 , splitterfromN68 , splitterfromN75 , splitterfromN8 , splitterN80ton149n76 , splitterN80ton64n76 , splitterN91ton93n345 , splitterN91ton262n345 , splitterN96ton90n360 , splitterN96ton273n360 , splitterfromn61 , splitterfromn63 , splittern65ton72N390 , splittern67ton160n69 , splitterfromn68 , splitterfromn70 , splitterfromn71 , splitterfromn73 , splitterfromn75 , splitterfromn78 , splittern81ton145N447 , splittern83ton179n88 , splitterfromn86 , splitterfromn92 , splitterfromn95 , splitterfromn98 , splitterfromn101 , splitterfromn104 , splitterfromn107 , splitterfromn110 , splitterfromn113 , splitterfromn119 , splitterfromn122 , splitterfromn125 , splitterfromn128 , splitterfromn131 , splitterfromn134 , splitterfromn137 , splitterfromn140 , splitterfromn144 , splitterfromn145 , splittern147ton148n208 , splitterfromn150 , splittern152ton164n210 , splittern162ton163n262 , splittern162ton207n262 , splittern162ton273n262 , splittern165ton166n175 , splitterfromn166 , splittern167ton168n201 , splittern168ton169n173 , splittern179ton253n346 , splittern179ton315n346 , splittern179ton221n346 , splittern192ton235n194 , splittern192ton193n194 , splittern193ton228n206 , splitterfromn194 , splittern198ton199n252 , splittern199ton245n204 , splitterfromn200 , splittern202ton203n247 , splittern204ton205n230 , splittern206ton214n297 , splittern210ton220n212 , splittern210ton211n212 , splittern211ton213n298 , splitterfromn212 , splittern213ton218n215 , splittern228ton229n233 , splittern245ton246n250 , splittern263ton264n282 , splittern266ton268n292 , splittern270ton329n272 , splittern270ton271n272 , splittern271ton328n306 , splitterfromn272 , splittern278ton344n280 , splittern278ton279n280 , splittern279ton343n304 , splittern279ton337n304 , splitterfromn280 , splittern286ton359n288 , splittern286ton287n288 , splittern287ton358n302 , splittern287ton352n302 , splitterfromn288 , splittern294ton314n296 , splittern294ton295n296 , splittern295ton313n300 , splitterfromn296 , splittern298ton299n312 , splittern300ton301n354 , splittern302ton303n339 , splittern304ton305n324 , splitterfromn307 , splittern322ton327n324 , splittern322ton323n324 , splittern337ton342n339 , splittern352ton357n354 ;

PI_AQFP N1_( clk_1 , N1 );
PI_AQFP N101_( clk_1 , N101 );
PI_AQFP N106_( clk_1 , N106 );
PI_AQFP N111_( clk_1 , N111 );
PI_AQFP N116_( clk_1 , N116 );
PI_AQFP N121_( clk_1 , N121 );
PI_AQFP N126_( clk_1 , N126 );
PI_AQFP N13_( clk_1 , N13 );
PI_AQFP N130_( clk_1 , N130 );
PI_AQFP N135_( clk_1 , N135 );
PI_AQFP N138_( clk_1 , N138 );
PI_AQFP N143_( clk_1 , N143 );
PI_AQFP N146_( clk_1 , N146 );
PI_AQFP N149_( clk_1 , N149 );
PI_AQFP N152_( clk_1 , N152 );
PI_AQFP N153_( clk_1 , N153 );
PI_AQFP N156_( clk_1 , N156 );
PI_AQFP N159_( clk_1 , N159 );
PI_AQFP N165_( clk_1 , N165 );
PI_AQFP N17_( clk_1 , N17 );
PI_AQFP N171_( clk_1 , N171 );
PI_AQFP N177_( clk_1 , N177 );
PI_AQFP N183_( clk_1 , N183 );
PI_AQFP N189_( clk_1 , N189 );
PI_AQFP N195_( clk_1 , N195 );
PI_AQFP N201_( clk_1 , N201 );
PI_AQFP N207_( clk_1 , N207 );
PI_AQFP N210_( clk_1 , N210 );
PI_AQFP N219_( clk_1 , N219 );
PI_AQFP N228_( clk_1 , N228 );
PI_AQFP N237_( clk_1 , N237 );
PI_AQFP N246_( clk_1 , N246 );
PI_AQFP N255_( clk_1 , N255 );
PI_AQFP N259_( clk_1 , N259 );
PI_AQFP N26_( clk_1 , N26 );
PI_AQFP N260_( clk_1 , N260 );
PI_AQFP N261_( clk_1 , N261 );
PI_AQFP N267_( clk_1 , N267 );
PI_AQFP N268_( clk_1 , N268 );
PI_AQFP N29_( clk_1 , N29 );
PI_AQFP N36_( clk_1 , N36 );
PI_AQFP N42_( clk_1 , N42 );
PI_AQFP N51_( clk_1 , N51 );
PI_AQFP N55_( clk_1 , N55 );
PI_AQFP N59_( clk_1 , N59 );
PI_AQFP N68_( clk_1 , N68 );
PI_AQFP N72_( clk_1 , N72 );
PI_AQFP N73_( clk_1 , N73 );
PI_AQFP N74_( clk_1 , N74 );
PI_AQFP N75_( clk_1 , N75 );
PI_AQFP N8_( clk_1 , N8 );
PI_AQFP N80_( clk_1 , N80 );
PI_AQFP N85_( clk_1 , N85 );
PI_AQFP N86_( clk_1 , N86 );
PI_AQFP N87_( clk_1 , N87 );
PI_AQFP N88_( clk_1 , N88 );
PI_AQFP N89_( clk_1 , N89 );
PI_AQFP N90_( clk_1 , N90 );
PI_AQFP N91_( clk_1 , N91 );
PI_AQFP N96_( clk_1 , N96 );
and_AQFP n61_( clk_4 , splitterN29ton61n84 , splitterfromN75 , 0 , 0 , n61 );
and_AQFP n62_( clk_1 , splitterN42ton62n77 , buf_splitterfromn61_n62_1 , 0 , 0 , n62 );
and_AQFP n63_( clk_5 , splitterN29ton61n84 , splitterfromN36 , 0 , 0 , n63 );
and_AQFP n64_( clk_2 , splitterN80ton64n76 , splitterfromn63 , 0 , 0 , n64 );
and_AQFP n65_( clk_2 , splitterN42ton62n77 , splitterfromn63 , 0 , 0 , n65 );
and_AQFP n66_( clk_3 , N85 , N86 , 0 , 0 , n66 );
and_AQFP n67_( clk_4 , splitterN1ton70n147 , splitterfromN8 , 0 , 0 , n67 );
and_AQFP n68_( clk_6 , buf_splitterfromN13_n68_1 , splitterN17ton68n283 , 0 , 0 , n68 );
and_AQFP n69_( clk_8 , buf_splittern67ton160n69_n69_1 , splitterfromn68 , 0 , 0 , n69 );
and_AQFP n70_( clk_3 , splitterN1ton70n147 , N26 , 0 , 0 , n70 );
and_AQFP n71_( clk_8 , splitterfromn68 , buf_splitterfromn70_n71_1 , 0 , 0 , n71 );
and_AQFP n72_( clk_8 , splittern65ton72N390 , splitterfromn71 , 1 , 0 , n72 );
and_AQFP n73_( clk_4 , splitterN59ton73n75 , splitterfromN75 , 0 , 0 , n73 );
and_AQFP n74_( clk_2 , splitterN80ton64n76 , buf_splitterfromn73_n74_1 , 0 , 0 , n74 );
and_AQFP n75_( clk_5 , splitterfromN36 , splitterN59ton73n75 , 0 , 0 , n75 );
and_AQFP n76_( clk_2 , splitterN80ton64n76 , splitterfromn75 , 0 , 0 , n76 );
and_AQFP n77_( clk_2 , splitterN42ton62n77 , splitterfromn75 , 0 , 0 , n77 );
or_AQFP n78_( clk_2 , N87 , N88 , 0 , 0 , n78 );
and_AQFP n79_( clk_4 , buf_N90_n79_1 , splitterfromn78 , 0 , 0 , n79 );
and_AQFP n80_( clk_8 , splittern65ton72N390 , splitterfromn71 , 0 , 0 , n80 );
and_AQFP n81_( clk_5 , splitterN51ton81n275 , splitterfromn70 , 0 , 0 , n81 );
and_AQFP n82_( clk_5 , splitterfromN13 , splitterN55ton82n263 , 0 , 0 , n82 );
and_AQFP n83_( clk_6 , splittern67ton160n69 , n82 , 0 , 0 , n83 );
and_AQFP n84_( clk_5 , splitterN29ton61n84 , splitterfromN68 , 0 , 0 , n84 );
and_AQFP n85_( clk_8 , splittern83ton179n88 , buf_n84_n85_1 , 0 , 0 , n85 );
and_AQFP n86_( clk_4 , splitterN59ton73n75 , splitterfromN68 , 0 , 0 , n86 );
and_AQFP n87_( clk_6 , buf_N74_n87_1 , splitterfromn86 , 0 , 0 , n87 );
and_AQFP n88_( clk_8 , splittern83ton179n88 , n87 , 0 , 0 , n88 );
and_AQFP n89_( clk_4 , buf_N89_n89_1 , splitterfromn78 , 0 , 0 , n89 );
or_AQFP n90_( clk_7 , splitterN130ton90n121 , splitterN96ton90n360 , 0 , 0 , n90 );
and_AQFP n91_( clk_7 , splitterN130ton90n121 , splitterN96ton90n360 , 0 , 0 , n91 );
and_AQFP n92_( clk_1 , n90 , n91 , 0 , 1 , n92 );
and_AQFP n93_( clk_5 , splitterN91ton93n345 , splitterfromn92 , 0 , 0 , n93 );
or_AQFP n94_( clk_5 , splitterN91ton93n345 , splitterfromn92 , 0 , 0 , n94 );
and_AQFP n95_( clk_7 , n93 , n94 , 1 , 0 , n95 );
or_AQFP n96_( clk_4 , splitterN121ton182n196 , splitterfromN135 , 0 , 0 , n96 );
and_AQFP n97_( clk_4 , splitterN121ton182n196 , splitterfromN135 , 0 , 0 , n97 );
and_AQFP n98_( clk_5 , n96 , n97 , 0 , 1 , n98 );
and_AQFP n99_( clk_8 , splitterN126ton100n163 , splitterfromn98 , 0 , 1 , n99 );
and_AQFP n100_( clk_8 , splitterN126ton100n163 , splitterfromn98 , 1 , 0 , n100 );
or_AQFP n101_( clk_1 , n99 , n100 , 0 , 0 , n101 );
and_AQFP n102_( clk_5 , splitterN101ton102n316 , splitterN106ton102n222 , 0 , 1 , n102 );
and_AQFP n103_( clk_5 , splitterN101ton102n316 , splitterN106ton102n222 , 1 , 0 , n103 );
or_AQFP n104_( clk_6 , n102 , n103 , 0 , 0 , n104 );
or_AQFP n105_( clk_5 , splitterN111ton105n207 , splitterN116ton105n190 , 0 , 0 , n105 );
and_AQFP n106_( clk_5 , splitterN111ton105n207 , splitterN116ton105n190 , 0 , 0 , n106 );
and_AQFP n107_( clk_6 , n105 , n106 , 0 , 1 , n107 );
or_AQFP n108_( clk_8 , splitterfromn104 , splitterfromn107 , 0 , 0 , n108 );
and_AQFP n109_( clk_8 , splitterfromn104 , splitterfromn107 , 0 , 0 , n109 );
and_AQFP n110_( clk_1 , n108 , n109 , 0 , 1 , n110 );
or_AQFP n111_( clk_5 , splitterfromn101 , splitterfromn110 , 0 , 0 , n111 );
and_AQFP n112_( clk_5 , splitterfromn101 , splitterfromn110 , 0 , 0 , n112 );
and_AQFP n113_( clk_7 , n111 , n112 , 0 , 1 , n113 );
and_AQFP n114_( clk_3 , splitterfromn95 , splitterfromn113 , 1 , 0 , n114 );
and_AQFP n115_( clk_3 , splitterfromn95 , splitterfromn113 , 0 , 1 , n115 );
or_AQFP n116_( clk_5 , n114 , n115 , 0 , 0 , n116 );
or_AQFP n117_( clk_4 , splitterN159ton117n272 , splitterN177ton117n296 , 0 , 0 , n117 );
and_AQFP n118_( clk_4 , splitterN159ton117n272 , splitterN177ton117n296 , 0 , 0 , n118 );
and_AQFP n119_( clk_5 , n117 , n118 , 0 , 1 , n119 );
and_AQFP n120_( clk_1 , splitterN130ton120n121 , splitterfromn119 , 0 , 1 , n120 );
and_AQFP n121_( clk_1 , splitterN130ton120n121 , splitterfromn119 , 1 , 0 , n121 );
or_AQFP n122_( clk_3 , n120 , n121 , 0 , 0 , n122 );
or_AQFP n123_( clk_4 , splitterN189ton123n194 , splitterN195ton123n200 , 0 , 0 , n123 );
and_AQFP n124_( clk_4 , splitterN189ton123n194 , splitterN195ton123n200 , 0 , 0 , n124 );
and_AQFP n125_( clk_5 , n123 , n124 , 0 , 1 , n125 );
and_AQFP n126_( clk_7 , splitterfromN207 , splitterfromn125 , 0 , 1 , n126 );
and_AQFP n127_( clk_7 , splitterfromN207 , splitterfromn125 , 1 , 0 , n127 );
or_AQFP n128_( clk_8 , n126 , n127 , 0 , 0 , n128 );
and_AQFP n129_( clk_4 , splitterN165ton129n280 , splitterN201ton129n167 , 1 , 0 , n129 );
and_AQFP n130_( clk_4 , splitterN165ton129n280 , splitterN201ton129n167 , 0 , 1 , n130 );
or_AQFP n131_( clk_5 , n129 , n130 , 0 , 0 , n131 );
and_AQFP n132_( clk_4 , splitterN171ton132n288 , splitterN183ton132n212 , 0 , 1 , n132 );
and_AQFP n133_( clk_4 , splitterN171ton132n288 , splitterN183ton132n212 , 1 , 0 , n133 );
or_AQFP n134_( clk_5 , n132 , n133 , 0 , 0 , n134 );
and_AQFP n135_( clk_7 , splitterfromn131 , splitterfromn134 , 0 , 1 , n135 );
and_AQFP n136_( clk_7 , splitterfromn131 , splitterfromn134 , 1 , 0 , n136 );
or_AQFP n137_( clk_8 , n135 , n136 , 0 , 0 , n137 );
and_AQFP n138_( clk_3 , splitterfromn128 , splitterfromn137 , 1 , 0 , n138 );
and_AQFP n139_( clk_2 , splitterfromn128 , splitterfromn137 , 0 , 1 , n139 );
or_AQFP n140_( clk_4 , n138 , n139 , 0 , 0 , n140 );
and_AQFP n141_( clk_7 , splitterfromn122 , splitterfromn140 , 0 , 1 , n141 );
and_AQFP n142_( clk_7 , splitterfromn122 , splitterfromn140 , 1 , 0 , n142 );
or_AQFP n143_( clk_1 , n141 , n142 , 0 , 0 , n143 );
and_AQFP n144_( clk_3 , N156 , splitterN59ton144n75 , 0 , 0 , n144 );
and_AQFP n145_( clk_7 , splittern81ton145N447 , splitterfromn144 , 0 , 1 , n145 );
and_AQFP n146_( clk_1 , splitterN17ton146n283 , splitterfromn145 , 0 , 0 , n146 );
and_AQFP n147_( clk_2 , buf_splitterN1ton70n147_n147_1 , n146 , 0 , 1 , n147 );
and_AQFP n148_( clk_4 , splitterfromN153 , splittern147ton148n208 , 0 , 1 , n148 );
and_AQFP n149_( clk_6 , splitterN80ton149n76 , splitterfromn61 , 0 , 0 , n149 );
and_AQFP n150_( clk_7 , splittern81ton145N447 , n149 , 0 , 0 , n150 );
and_AQFP n151_( clk_1 , splitterN55ton151n263 , splitterfromn150 , 0 , 0 , n151 );
and_AQFP n152_( clk_2 , splitterN268ton152n331 , n151 , 1 , 0 , n152 );
and_AQFP n153_( clk_5 , splitterN17ton153n283 , splitterN42ton153n77 , 0 , 1 , n153 );
and_AQFP n154_( clk_5 , splitterN17ton153n283 , splitterN42ton153n77 , 1 , 0 , n154 );
or_AQFP n155_( clk_6 , n153 , n154 , 0 , 0 , n155 );
and_AQFP n156_( clk_7 , splittern81ton145N447 , splitterfromn144 , 0 , 0 , n156 );
and_AQFP n157_( clk_8 , n155 , n156 , 0 , 0 , n157 );
and_AQFP n158_( clk_7 , splitterN42ton158n77 , splitterfromn73 , 0 , 0 , n158 );
and_AQFP n159_( clk_5 , splitterN17ton153n283 , splitterN51ton159n275 , 0 , 0 , n159 );
and_AQFP n160_( clk_6 , splittern67ton160n69 , n159 , 0 , 0 , n160 );
and_AQFP n161_( clk_8 , n158 , n160 , 1 , 0 , n161 );
or_AQFP n162_( clk_1 , n157 , n161 , 0 , 0 , n162 );
and_AQFP n163_( clk_3 , buf_splitterN126ton100n163_n163_1 , splittern162ton163n262 , 0 , 0 , n163 );
or_AQFP n164_( clk_4 , splittern152ton164n210 , n163 , 0 , 0 , n164 );
or_AQFP n165_( clk_5 , n148 , n164 , 0 , 0 , n165 );
or_AQFP n166_( clk_7 , splitterN201ton166n167 , splittern165ton166n175 , 0 , 0 , n166 );
and_AQFP n167_( clk_7 , splitterN201ton166n167 , splittern165ton166n175 , 0 , 0 , n167 );
and_AQFP n168_( clk_1 , splitterfromn166 , splittern167ton168n201 , 0 , 1 , n168 );
and_AQFP n169_( clk_3 , splitterN261ton169n170 , splittern168ton169n173 , 0 , 0 , n169 );
or_AQFP n170_( clk_3 , splitterN261ton169n170 , splittern168ton169n173 , 0 , 0 , n170 );
and_AQFP n171_( clk_4 , splitterN219ton171n325 , n170 , 0 , 0 , n171 );
and_AQFP n172_( clk_5 , n169 , n171 , 1 , 0 , n172 );
and_AQFP n173_( clk_3 , splitterN228ton173n342 , splittern168ton169n173 , 0 , 0 , n173 );
and_AQFP n174_( clk_1 , splitterN237ton174n328 , splittern167ton168n201 , 0 , 0 , n174 );
and_AQFP n175_( clk_7 , splitterN246ton175n359 , splittern165ton166n175 , 0 , 0 , n175 );
and_AQFP n176_( clk_3 , splitterN42ton176n77 , N72 , 0 , 0 , n176 );
and_AQFP n177_( clk_4 , buf_N73_n177_1 , n176 , 0 , 0 , n177 );
and_AQFP n178_( clk_6 , splitterfromn86 , n177 , 0 , 0 , n178 );
and_AQFP n179_( clk_8 , splittern83ton179n88 , n178 , 0 , 0 , n179 );
and_AQFP n180_( clk_2 , splitterN201ton180n167 , splittern179ton253n346 , 0 , 0 , n180 );
and_AQFP n181_( clk_3 , splitterN255ton181n254 , N267 , 0 , 0 , n181 );
and_AQFP n182_( clk_4 , splitterN121ton182n196 , splitterN210ton182n345 , 0 , 0 , n182 );
or_AQFP n183_( clk_6 , buf_n181_n183_1 , n182 , 0 , 0 , n183 );
or_AQFP n184_( clk_3 , n180 , buf_n183_n184_1 , 0 , 0 , n184 );
or_AQFP n185_( clk_8 , n175 , buf_n184_n185_1 , 0 , 0 , n185 );
or_AQFP n186_( clk_2 , n174 , n185 , 0 , 0 , n186 );
or_AQFP n187_( clk_4 , n173 , n186 , 0 , 0 , n187 );
or_AQFP n188_( clk_6 , n172 , n187 , 0 , 0 , n188 );
and_AQFP n189_( clk_4 , buf_splitterfromN146_n189_1 , splittern147ton148n208 , 0 , 1 , n189 );
and_AQFP n190_( clk_3 , buf_splitterN116ton105n190_n190_1 , splittern162ton163n262 , 0 , 0 , n190 );
or_AQFP n191_( clk_5 , splittern152ton164n210 , n190 , 0 , 0 , n191 );
or_AQFP n192_( clk_6 , n189 , n191 , 0 , 0 , n192 );
and_AQFP n193_( clk_3 , splitterN189ton193n194 , splittern192ton193n194 , 0 , 0 , n193 );
or_AQFP n194_( clk_3 , splitterN189ton193n194 , splittern192ton193n194 , 0 , 0 , n194 );
and_AQFP n195_( clk_4 , splitterfromN149 , splittern147ton148n208 , 0 , 1 , n195 );
and_AQFP n196_( clk_3 , buf_splitterN121ton182n196_n196_1 , splittern162ton163n262 , 0 , 0 , n196 );
or_AQFP n197_( clk_4 , splittern152ton164n210 , n196 , 0 , 0 , n197 );
or_AQFP n198_( clk_5 , n195 , n197 , 0 , 0 , n198 );
and_AQFP n199_( clk_8 , splitterN195ton199n200 , splittern198ton199n252 , 0 , 0 , n199 );
or_AQFP n200_( clk_8 , splitterN195ton199n200 , splittern198ton199n252 , 0 , 0 , n200 );
or_AQFP n201_( clk_1 , splitterN261ton201n170 , splittern167ton168n201 , 0 , 0 , n201 );
and_AQFP n202_( clk_2 , splitterfromn166 , n201 , 0 , 0 , n202 );
and_AQFP n203_( clk_4 , splitterfromn200 , splittern202ton203n247 , 0 , 0 , n203 );
or_AQFP n204_( clk_5 , buf_splittern199ton245n204_n204_1 , n203 , 0 , 0 , n204 );
and_AQFP n205_( clk_7 , splitterfromn194 , splittern204ton205n230 , 0 , 0 , n205 );
or_AQFP n206_( clk_8 , buf_splittern193ton228n206_n206_1 , n205 , 0 , 0 , n206 );
and_AQFP n207_( clk_4 , buf_splitterN111ton105n207_n207_1 , splittern162ton207n262 , 0 , 0 , n207 );
and_AQFP n208_( clk_4 , splitterfromN143 , splittern147ton148n208 , 0 , 1 , n208 );
or_AQFP n209_( clk_5 , n207 , n208 , 0 , 0 , n209 );
or_AQFP n210_( clk_6 , buf_splittern152ton164n210_n210_1 , n209 , 0 , 0 , n210 );
and_AQFP n211_( clk_4 , splitterN183ton211n212 , splittern210ton211n212 , 0 , 0 , n211 );
or_AQFP n212_( clk_4 , splitterN183ton211n212 , splittern210ton211n212 , 0 , 0 , n212 );
and_AQFP n213_( clk_7 , splittern211ton213n298 , splitterfromn212 , 1 , 0 , n213 );
or_AQFP n214_( clk_2 , splittern206ton214n297 , splittern213ton218n215 , 0 , 0 , n214 );
and_AQFP n215_( clk_2 , splittern206ton214n297 , splittern213ton218n215 , 0 , 0 , n215 );
and_AQFP n216_( clk_3 , n214 , n215 , 0 , 1 , n216 );
and_AQFP n217_( clk_5 , splitterN219ton217n325 , n216 , 0 , 0 , n217 );
and_AQFP n218_( clk_1 , splitterN228ton218n342 , splittern213ton218n215 , 0 , 0 , n218 );
and_AQFP n219_( clk_7 , splitterN237ton219n328 , splittern211ton213n298 , 0 , 0 , n219 );
and_AQFP n220_( clk_1 , splitterN246ton235n359 , splittern210ton220n212 , 0 , 0 , n220 );
and_AQFP n221_( clk_6 , splitterN183ton221n212 , splittern179ton221n346 , 0 , 0 , n221 );
and_AQFP n222_( clk_6 , buf_splitterN106ton289n222_n222_1 , splitterN210ton222n345 , 0 , 0 , n222 );
or_AQFP n223_( clk_8 , n221 , n222 , 0 , 0 , n223 );
or_AQFP n224_( clk_2 , n220 , n223 , 0 , 0 , n224 );
or_AQFP n225_( clk_8 , n219 , buf_n224_n225_1 , 0 , 0 , n225 );
or_AQFP n226_( clk_2 , n218 , n225 , 0 , 0 , n226 );
or_AQFP n227_( clk_6 , n217 , buf_n226_n227_1 , 0 , 0 , n227 );
and_AQFP n228_( clk_6 , splittern193ton228n206 , splitterfromn194 , 1 , 0 , n228 );
or_AQFP n229_( clk_8 , splittern204ton205n230 , splittern228ton229n233 , 0 , 0 , n229 );
and_AQFP n230_( clk_8 , splittern204ton205n230 , splittern228ton229n233 , 0 , 0 , n230 );
and_AQFP n231_( clk_1 , n229 , n230 , 0 , 1 , n231 );
and_AQFP n232_( clk_2 , splitterN219ton232n325 , n231 , 0 , 0 , n232 );
and_AQFP n233_( clk_8 , splitterN228ton233n342 , splittern228ton229n233 , 0 , 0 , n233 );
and_AQFP n234_( clk_6 , splitterN237ton234n328 , splittern193ton228n206 , 0 , 0 , n234 );
and_AQFP n235_( clk_8 , splitterN246ton235n359 , splittern192ton235n194 , 0 , 0 , n235 );
and_AQFP n236_( clk_2 , splitterN189ton236n194 , splittern179ton253n346 , 0 , 0 , n236 );
and_AQFP n237_( clk_5 , splitterN111ton105n207 , splitterN210ton182n345 , 0 , 0 , n237 );
and_AQFP n238_( clk_3 , splitterN255ton181n254 , N259 , 0 , 0 , n238 );
or_AQFP n239_( clk_6 , n237 , buf_n238_n239_1 , 0 , 0 , n239 );
or_AQFP n240_( clk_3 , n236 , buf_n239_n240_1 , 0 , 0 , n240 );
or_AQFP n241_( clk_1 , n235 , buf_n240_n241_1 , 0 , 0 , n241 );
or_AQFP n242_( clk_7 , n234 , buf_n241_n242_1 , 0 , 0 , n242 );
or_AQFP n243_( clk_1 , n233 , n242 , 0 , 0 , n243 );
or_AQFP n244_( clk_4 , n232 , buf_n243_n244_1 , 0 , 0 , n244 );
and_AQFP n245_( clk_3 , splittern199ton245n204 , splitterfromn200 , 1 , 0 , n245 );
or_AQFP n246_( clk_5 , splittern202ton203n247 , splittern245ton246n250 , 0 , 0 , n246 );
and_AQFP n247_( clk_5 , splittern202ton203n247 , splittern245ton246n250 , 0 , 0 , n247 );
and_AQFP n248_( clk_6 , n246 , n247 , 0 , 1 , n248 );
and_AQFP n249_( clk_7 , splitterN219ton249n325 , n248 , 0 , 0 , n249 );
and_AQFP n250_( clk_5 , splitterN228ton250n342 , splittern245ton246n250 , 0 , 0 , n250 );
and_AQFP n251_( clk_3 , splitterN237ton251n328 , splittern199ton245n204 , 0 , 0 , n251 );
and_AQFP n252_( clk_8 , splitterN246ton235n359 , splittern198ton199n252 , 0 , 0 , n252 );
and_AQFP n253_( clk_2 , splitterN195ton253n200 , splittern179ton253n346 , 0 , 0 , n253 );
and_AQFP n254_( clk_4 , splitterN255ton181n254 , buf_N260_n254_1 , 0 , 0 , n254 );
and_AQFP n255_( clk_5 , splitterN116ton105n190 , splitterN210ton182n345 , 0 , 0 , n255 );
or_AQFP n256_( clk_6 , n254 , n255 , 0 , 0 , n256 );
or_AQFP n257_( clk_3 , n253 , buf_n256_n257_1 , 0 , 0 , n257 );
or_AQFP n258_( clk_1 , n252 , buf_n257_n258_1 , 0 , 0 , n258 );
or_AQFP n259_( clk_4 , n251 , buf_n258_n259_1 , 0 , 0 , n259 );
or_AQFP n260_( clk_6 , n250 , n259 , 0 , 0 , n260 );
or_AQFP n261_( clk_1 , n249 , buf_n260_n261_1 , 0 , 0 , n261 );
and_AQFP n262_( clk_6 , splitterN91ton262n345 , splittern162ton273n262 , 0 , 0 , n262 );
and_AQFP n263_( clk_1 , splitterN55ton151n263 , splitterfromn145 , 0 , 0 , n263 );
and_AQFP n264_( clk_4 , splitterfromN143 , splittern263ton264n282 , 0 , 0 , n264 );
and_AQFP n265_( clk_7 , splitterN17ton68n283 , splitterN268ton265n331 , 0 , 1 , n265 );
and_AQFP n266_( clk_1 , splitterfromn150 , n265 , 0 , 0 , n266 );
and_AQFP n267_( clk_1 , splitterN138ton291n283 , buf_splitterfromN8_n267_1 , 0 , 0 , n267 );
or_AQFP n268_( clk_3 , splittern266ton268n292 , n267 , 0 , 0 , n268 );
or_AQFP n269_( clk_5 , n264 , n268 , 0 , 0 , n269 );
or_AQFP n270_( clk_7 , n262 , n269 , 0 , 0 , n270 );
and_AQFP n271_( clk_5 , splitterN159ton271n272 , splittern270ton271n272 , 0 , 0 , n271 );
or_AQFP n272_( clk_5 , splitterN159ton271n272 , splittern270ton271n272 , 0 , 0 , n272 );
and_AQFP n273_( clk_5 , splitterN96ton273n360 , splittern162ton273n262 , 0 , 0 , n273 );
and_AQFP n274_( clk_3 , splitterfromN146 , splittern263ton264n282 , 0 , 0 , n274 );
and_AQFP n275_( clk_1 , splitterN138ton291n283 , buf_splitterN51ton81n275_n275_1 , 0 , 0 , n275 );
or_AQFP n276_( clk_3 , splittern266ton268n292 , n275 , 0 , 0 , n276 );
or_AQFP n277_( clk_5 , n274 , n276 , 0 , 0 , n277 );
or_AQFP n278_( clk_7 , n273 , n277 , 0 , 0 , n278 );
and_AQFP n279_( clk_5 , splitterN165ton279n280 , splittern278ton279n280 , 0 , 0 , n279 );
or_AQFP n280_( clk_5 , splitterN165ton279n280 , splittern278ton279n280 , 0 , 0 , n280 );
and_AQFP n281_( clk_5 , splitterN101ton281n316 , splittern162ton273n262 , 0 , 0 , n281 );
and_AQFP n282_( clk_3 , splitterfromN149 , splittern263ton264n282 , 0 , 0 , n282 );
and_AQFP n283_( clk_1 , splitterN138ton291n283 , splitterN17ton146n283 , 0 , 0 , n283 );
or_AQFP n284_( clk_3 , splittern266ton268n292 , n283 , 0 , 0 , n284 );
or_AQFP n285_( clk_5 , n282 , n284 , 0 , 0 , n285 );
or_AQFP n286_( clk_7 , n281 , n285 , 0 , 0 , n286 );
and_AQFP n287_( clk_5 , splitterN171ton287n288 , splittern286ton287n288 , 0 , 0 , n287 );
or_AQFP n288_( clk_5 , splitterN171ton287n288 , splittern286ton287n288 , 0 , 0 , n288 );
and_AQFP n289_( clk_5 , splitterN106ton289n222 , splittern162ton273n262 , 0 , 0 , n289 );
and_AQFP n290_( clk_3 , splitterfromN153 , splittern263ton264n282 , 0 , 0 , n290 );
and_AQFP n291_( clk_8 , splitterN138ton291n283 , buf_N152_n291_1 , 0 , 0 , n291 );
or_AQFP n292_( clk_3 , splittern266ton268n292 , buf_n291_n292_1 , 0 , 0 , n292 );
or_AQFP n293_( clk_5 , n290 , n292 , 0 , 0 , n293 );
or_AQFP n294_( clk_7 , n289 , n293 , 0 , 0 , n294 );
and_AQFP n295_( clk_5 , splitterN177ton295n296 , splittern294ton295n296 , 0 , 0 , n295 );
or_AQFP n296_( clk_5 , splitterN177ton295n296 , splittern294ton295n296 , 0 , 0 , n296 );
and_AQFP n297_( clk_2 , splittern206ton214n297 , buf_splitterfromn212_n297_1 , 0 , 0 , n297 );
or_AQFP n298_( clk_3 , buf_splittern211ton213n298_n298_1 , n297 , 0 , 0 , n298 );
and_AQFP n299_( clk_5 , buf_splitterfromn296_n299_1 , splittern298ton299n312 , 0 , 0 , n299 );
or_AQFP n300_( clk_6 , buf_splittern295ton313n300_n300_1 , n299 , 0 , 0 , n300 );
and_AQFP n301_( clk_8 , buf_splitterfromn288_n301_1 , splittern300ton301n354 , 0 , 0 , n301 );
or_AQFP n302_( clk_1 , buf_splittern287ton352n302_n302_1 , n301 , 0 , 0 , n302 );
and_AQFP n303_( clk_3 , buf_splitterfromn280_n303_1 , splittern302ton303n339 , 0 , 0 , n303 );
or_AQFP n304_( clk_4 , buf_splittern279ton337n304_n304_1 , n303 , 0 , 0 , n304 );
and_AQFP n305_( clk_6 , buf_splitterfromn272_n305_1 , splittern304ton305n324 , 0 , 0 , n305 );
or_AQFP n306_( clk_7 , buf_splittern271ton328n306_n306_1 , n305 , 0 , 0 , n306 );
and_AQFP n307_( clk_2 , splittern295ton313n300 , splitterfromn296 , 1 , 0 , n307 );
and_AQFP n308_( clk_5 , splitterN219ton217n325 , splittern298ton299n312 , 0 , 1 , n308 );
or_AQFP n309_( clk_6 , splitterN228ton309n342 , n308 , 0 , 0 , n309 );
and_AQFP n310_( clk_7 , buf_splitterfromn307_n310_1 , n309 , 0 , 0 , n310 );
and_AQFP n311_( clk_5 , splitterN219ton217n325 , splitterfromn307 , 0 , 1 , n311 );
and_AQFP n312_( clk_6 , splittern298ton299n312 , n311 , 0 , 0 , n312 );
and_AQFP n313_( clk_2 , splitterN237ton313n328 , splittern295ton313n300 , 0 , 0 , n313 );
and_AQFP n314_( clk_2 , splitterN246ton314n359 , splittern294ton314n296 , 0 , 0 , n314 );
and_AQFP n315_( clk_5 , splitterN177ton315n296 , splittern179ton315n346 , 0 , 0 , n315 );
and_AQFP n316_( clk_5 , splitterN101ton281n316 , splitterN210ton316n345 , 0 , 0 , n316 );
or_AQFP n317_( clk_7 , n315 , n316 , 0 , 0 , n317 );
or_AQFP n318_( clk_3 , n314 , buf_n317_n318_1 , 0 , 0 , n318 );
or_AQFP n319_( clk_4 , n313 , buf_n318_n319_1 , 0 , 0 , n319 );
or_AQFP n320_( clk_7 , n312 , buf_n319_n320_1 , 0 , 0 , n320 );
or_AQFP n321_( clk_1 , n310 , n320 , 0 , 0 , n321 );
and_AQFP n322_( clk_7 , splittern271ton328n306 , splitterfromn272 , 1 , 0 , n322 );
or_AQFP n323_( clk_6 , splittern304ton305n324 , splittern322ton323n324 , 0 , 0 , n323 );
and_AQFP n324_( clk_6 , splittern304ton305n324 , splittern322ton323n324 , 0 , 0 , n324 );
and_AQFP n325_( clk_7 , buf_splitterN219ton340n325_n325_1 , n324 , 0 , 1 , n325 );
and_AQFP n326_( clk_8 , n323 , n325 , 0 , 0 , n326 );
and_AQFP n327_( clk_2 , splitterN228ton327n342 , splittern322ton327n324 , 0 , 0 , n327 );
and_AQFP n328_( clk_6 , splitterN237ton343n328 , splittern271ton328n306 , 0 , 0 , n328 );
and_AQFP n329_( clk_2 , splitterN246ton314n359 , splittern270ton329n272 , 0 , 0 , n329 );
and_AQFP n330_( clk_6 , splitterN159ton330n272 , splittern179ton221n346 , 0 , 0 , n330 );
and_AQFP n331_( clk_6 , splitterN210ton222n345 , buf_splitterN268ton152n331_n331_1 , 0 , 0 , n331 );
or_AQFP n332_( clk_8 , n330 , n331 , 0 , 0 , n332 );
or_AQFP n333_( clk_3 , n329 , buf_n332_n333_1 , 0 , 0 , n333 );
or_AQFP n334_( clk_7 , n328 , buf_n333_n334_1 , 0 , 0 , n334 );
or_AQFP n335_( clk_3 , n327 , buf_n334_n335_1 , 0 , 0 , n335 );
or_AQFP n336_( clk_1 , n326 , buf_n335_n336_1 , 0 , 0 , n336 );
and_AQFP n337_( clk_7 , splittern279ton337n304 , splitterfromn280 , 1 , 0 , n337 );
and_AQFP n338_( clk_3 , splittern302ton303n339 , splittern337ton342n339 , 0 , 0 , n338 );
or_AQFP n339_( clk_3 , splittern302ton303n339 , splittern337ton342n339 , 0 , 0 , n339 );
and_AQFP n340_( clk_4 , splitterN219ton340n325 , n339 , 0 , 0 , n340 );
and_AQFP n341_( clk_5 , n338 , n340 , 1 , 0 , n341 );
and_AQFP n342_( clk_2 , splitterN228ton327n342 , splittern337ton342n339 , 0 , 0 , n342 );
and_AQFP n343_( clk_5 , splitterN237ton343n328 , splittern279ton343n304 , 0 , 0 , n343 );
and_AQFP n344_( clk_2 , splitterN246ton314n359 , splittern278ton344n280 , 0 , 0 , n344 );
and_AQFP n345_( clk_7 , splitterN210ton222n345 , splitterN91ton262n345 , 0 , 0 , n345 );
and_AQFP n346_( clk_7 , splitterN165ton346n280 , splittern179ton221n346 , 0 , 0 , n346 );
or_AQFP n347_( clk_1 , n345 , n346 , 0 , 0 , n347 );
or_AQFP n348_( clk_3 , n344 , n347 , 0 , 0 , n348 );
or_AQFP n349_( clk_6 , n343 , buf_n348_n349_1 , 0 , 0 , n349 );
or_AQFP n350_( clk_3 , n342 , buf_n349_n350_1 , 0 , 0 , n350 );
or_AQFP n351_( clk_6 , n341 , buf_n350_n351_1 , 0 , 0 , n351 );
and_AQFP n352_( clk_4 , splittern287ton352n302 , splitterfromn288 , 1 , 0 , n352 );
and_AQFP n353_( clk_8 , splittern300ton301n354 , splittern352ton357n354 , 0 , 0 , n353 );
or_AQFP n354_( clk_8 , splittern300ton301n354 , splittern352ton357n354 , 0 , 0 , n354 );
and_AQFP n355_( clk_1 , splitterN219ton355n325 , n354 , 0 , 0 , n355 );
and_AQFP n356_( clk_2 , n353 , n355 , 1 , 0 , n356 );
and_AQFP n357_( clk_7 , splitterN228ton357n342 , splittern352ton357n354 , 0 , 0 , n357 );
and_AQFP n358_( clk_3 , splitterN237ton358n328 , splittern287ton358n302 , 0 , 0 , n358 );
and_AQFP n359_( clk_2 , splitterN246ton314n359 , splittern286ton359n288 , 0 , 0 , n359 );
and_AQFP n360_( clk_6 , splitterN210ton222n345 , buf_splitterN96ton273n360_n360_1 , 0 , 0 , n360 );
and_AQFP n361_( clk_6 , splitterN171ton361n288 , splittern179ton221n346 , 0 , 0 , n361 );
or_AQFP n362_( clk_8 , n360 , n361 , 0 , 0 , n362 );
or_AQFP n363_( clk_3 , n359 , buf_n362_n363_1 , 0 , 0 , n363 );
or_AQFP n364_( clk_4 , n358 , buf_n363_n364_1 , 0 , 0 , n364 );
or_AQFP n365_( clk_8 , n357 , buf_n364_n365_1 , 0 , 0 , n365 );
or_AQFP n366_( clk_3 , n356 , buf_n365_n366_1 , 0 , 0 , n366 );
PO_AQFP N388_( clk_2 , buf_n62_N388_1 , 0 , N388 );
PO_AQFP N389_( clk_2 , buf_n64_N389_1 , 0 , N389 );
PO_AQFP N390_( clk_2 , buf_splittern65ton72N390_N390_1 , 0 , N390 );
PO_AQFP N391_( clk_2 , buf_n66_N391_1 , 0 , N391 );
PO_AQFP N418_( clk_2 , buf_n69_N418_1 , 0 , N418 );
PO_AQFP N419_( clk_2 , n72 , 1 , N419 );
PO_AQFP N420_( clk_2 , buf_n74_N420_1 , 1 , N420 );
PO_AQFP N421_( clk_2 , buf_n76_N421_1 , 1 , N421 );
PO_AQFP N422_( clk_2 , buf_n77_N422_1 , 1 , N422 );
PO_AQFP N423_( clk_2 , buf_n79_N423_1 , 0 , N423 );
PO_AQFP N446_( clk_2 , n80 , 1 , N446 );
PO_AQFP N447_( clk_2 , buf_splittern81ton145N447_N447_1 , 0 , N447 );
PO_AQFP N448_( clk_2 , buf_n85_N448_1 , 0 , N448 );
PO_AQFP N449_( clk_2 , buf_n88_N449_1 , 0 , N449 );
PO_AQFP N450_( clk_2 , buf_n89_N450_1 , 0 , N450 );
PO_AQFP N767_( clk_2 , buf_n116_N767_1 , 0 , N767 );
PO_AQFP N768_( clk_2 , buf_n143_N768_1 , 0 , N768 );
PO_AQFP N850_( clk_2 , buf_n188_N850_1 , 0 , N850 );
PO_AQFP N863_( clk_2 , buf_n227_N863_1 , 0 , N863 );
PO_AQFP N864_( clk_2 , buf_n244_N864_1 , 0 , N864 );
PO_AQFP N865_( clk_2 , buf_n261_N865_1 , 0 , N865 );
PO_AQFP N866_( clk_2 , buf_n306_N866_1 , 0 , N866 );
PO_AQFP N874_( clk_2 , buf_n321_N874_1 , 0 , N874 );
PO_AQFP N878_( clk_2 , n336 , 0 , N878 );
PO_AQFP N879_( clk_2 , buf_n351_N879_1 , 0 , N879 );
PO_AQFP N880_( clk_2 , buf_n366_N880_1 , 0 , N880 );
buf_AQFP buf_N101_splitterN101ton102n316_1_( clk_3 , N101 , 0 , buf_N101_splitterN101ton102n316_1 );
buf_AQFP buf_N111_splitterN111ton105n207_1_( clk_3 , N111 , 0 , buf_N111_splitterN111ton105n207_1 );
buf_AQFP buf_N116_splitterN116ton105n190_1_( clk_3 , N116 , 0 , buf_N116_splitterN116ton105n190_1 );
buf_AQFP buf_N126_splitterN126ton100n163_2_( clk_3 , N126 , 0 , buf_N126_splitterN126ton100n163_2 );
buf_AQFP buf_N126_splitterN126ton100n163_1_( clk_5 , buf_N126_splitterN126ton100n163_2 , 0 , buf_N126_splitterN126ton100n163_1 );
buf_AQFP buf_N130_splitterN130ton90n121_1_( clk_3 , N130 , 0 , buf_N130_splitterN130ton90n121_1 );
buf_AQFP buf_N138_splitterN138ton291n283_2_( clk_3 , N138 , 0 , buf_N138_splitterN138ton291n283_2 );
buf_AQFP buf_N138_splitterN138ton291n283_1_( clk_5 , buf_N138_splitterN138ton291n283_2 , 0 , buf_N138_splitterN138ton291n283_1 );
buf_AQFP buf_N143_splitterfromN143_4_( clk_3 , N143 , 0 , buf_N143_splitterfromN143_4 );
buf_AQFP buf_N143_splitterfromN143_3_( clk_5 , buf_N143_splitterfromN143_4 , 0 , buf_N143_splitterfromN143_3 );
buf_AQFP buf_N143_splitterfromN143_2_( clk_7 , buf_N143_splitterfromN143_3 , 0 , buf_N143_splitterfromN143_2 );
buf_AQFP buf_N143_splitterfromN143_1_( clk_1 , buf_N143_splitterfromN143_2 , 0 , buf_N143_splitterfromN143_1 );
buf_AQFP buf_N146_splitterfromN146_3_( clk_3 , N146 , 0 , buf_N146_splitterfromN146_3 );
buf_AQFP buf_N146_splitterfromN146_2_( clk_5 , buf_N146_splitterfromN146_3 , 0 , buf_N146_splitterfromN146_2 );
buf_AQFP buf_N146_splitterfromN146_1_( clk_7 , buf_N146_splitterfromN146_2 , 0 , buf_N146_splitterfromN146_1 );
buf_AQFP buf_N149_splitterfromN149_4_( clk_3 , N149 , 0 , buf_N149_splitterfromN149_4 );
buf_AQFP buf_N149_splitterfromN149_3_( clk_5 , buf_N149_splitterfromN149_4 , 0 , buf_N149_splitterfromN149_3 );
buf_AQFP buf_N149_splitterfromN149_2_( clk_7 , buf_N149_splitterfromN149_3 , 0 , buf_N149_splitterfromN149_2 );
buf_AQFP buf_N149_splitterfromN149_1_( clk_1 , buf_N149_splitterfromN149_2 , 0 , buf_N149_splitterfromN149_1 );
buf_AQFP buf_N152_n291_3_( clk_3 , N152 , 0 , buf_N152_n291_3 );
buf_AQFP buf_N152_n291_2_( clk_5 , buf_N152_n291_3 , 0 , buf_N152_n291_2 );
buf_AQFP buf_N152_n291_1_( clk_7 , buf_N152_n291_2 , 0 , buf_N152_n291_1 );
buf_AQFP buf_N153_splitterfromN153_4_( clk_3 , N153 , 0 , buf_N153_splitterfromN153_4 );
buf_AQFP buf_N153_splitterfromN153_3_( clk_5 , buf_N153_splitterfromN153_4 , 0 , buf_N153_splitterfromN153_3 );
buf_AQFP buf_N153_splitterfromN153_2_( clk_7 , buf_N153_splitterfromN153_3 , 0 , buf_N153_splitterfromN153_2 );
buf_AQFP buf_N153_splitterfromN153_1_( clk_1 , buf_N153_splitterfromN153_2 , 0 , buf_N153_splitterfromN153_1 );
buf_AQFP buf_N207_splitterfromN207_1_( clk_3 , N207 , 0 , buf_N207_splitterfromN207_1 );
buf_AQFP buf_N219_splitterN219ton171n325_8_( clk_3 , N219 , 0 , buf_N219_splitterN219ton171n325_8 );
buf_AQFP buf_N219_splitterN219ton171n325_7_( clk_5 , buf_N219_splitterN219ton171n325_8 , 0 , buf_N219_splitterN219ton171n325_7 );
buf_AQFP buf_N219_splitterN219ton171n325_6_( clk_7 , buf_N219_splitterN219ton171n325_7 , 0 , buf_N219_splitterN219ton171n325_6 );
buf_AQFP buf_N219_splitterN219ton171n325_5_( clk_1 , buf_N219_splitterN219ton171n325_6 , 0 , buf_N219_splitterN219ton171n325_5 );
buf_AQFP buf_N219_splitterN219ton171n325_4_( clk_3 , buf_N219_splitterN219ton171n325_5 , 0 , buf_N219_splitterN219ton171n325_4 );
buf_AQFP buf_N219_splitterN219ton171n325_3_( clk_5 , buf_N219_splitterN219ton171n325_4 , 0 , buf_N219_splitterN219ton171n325_3 );
buf_AQFP buf_N219_splitterN219ton171n325_2_( clk_7 , buf_N219_splitterN219ton171n325_3 , 0 , buf_N219_splitterN219ton171n325_2 );
buf_AQFP buf_N219_splitterN219ton171n325_1_( clk_1 , buf_N219_splitterN219ton171n325_2 , 0 , buf_N219_splitterN219ton171n325_1 );
buf_AQFP buf_N228_splitterN228ton173n342_7_( clk_3 , N228 , 0 , buf_N228_splitterN228ton173n342_7 );
buf_AQFP buf_N228_splitterN228ton173n342_6_( clk_5 , buf_N228_splitterN228ton173n342_7 , 0 , buf_N228_splitterN228ton173n342_6 );
buf_AQFP buf_N228_splitterN228ton173n342_5_( clk_7 , buf_N228_splitterN228ton173n342_6 , 0 , buf_N228_splitterN228ton173n342_5 );
buf_AQFP buf_N228_splitterN228ton173n342_4_( clk_1 , buf_N228_splitterN228ton173n342_5 , 0 , buf_N228_splitterN228ton173n342_4 );
buf_AQFP buf_N228_splitterN228ton173n342_3_( clk_3 , buf_N228_splitterN228ton173n342_4 , 0 , buf_N228_splitterN228ton173n342_3 );
buf_AQFP buf_N228_splitterN228ton173n342_2_( clk_5 , buf_N228_splitterN228ton173n342_3 , 0 , buf_N228_splitterN228ton173n342_2 );
buf_AQFP buf_N228_splitterN228ton173n342_1_( clk_7 , buf_N228_splitterN228ton173n342_2 , 0 , buf_N228_splitterN228ton173n342_1 );
buf_AQFP buf_N237_splitterN237ton174n328_6_( clk_3 , N237 , 0 , buf_N237_splitterN237ton174n328_6 );
buf_AQFP buf_N237_splitterN237ton174n328_5_( clk_5 , buf_N237_splitterN237ton174n328_6 , 0 , buf_N237_splitterN237ton174n328_5 );
buf_AQFP buf_N237_splitterN237ton174n328_4_( clk_7 , buf_N237_splitterN237ton174n328_5 , 0 , buf_N237_splitterN237ton174n328_4 );
buf_AQFP buf_N237_splitterN237ton174n328_3_( clk_1 , buf_N237_splitterN237ton174n328_4 , 0 , buf_N237_splitterN237ton174n328_3 );
buf_AQFP buf_N237_splitterN237ton174n328_2_( clk_3 , buf_N237_splitterN237ton174n328_3 , 0 , buf_N237_splitterN237ton174n328_2 );
buf_AQFP buf_N237_splitterN237ton174n328_1_( clk_5 , buf_N237_splitterN237ton174n328_2 , 0 , buf_N237_splitterN237ton174n328_1 );
buf_AQFP buf_N246_splitterN246ton175n359_5_( clk_3 , N246 , 0 , buf_N246_splitterN246ton175n359_5 );
buf_AQFP buf_N246_splitterN246ton175n359_4_( clk_5 , buf_N246_splitterN246ton175n359_5 , 0 , buf_N246_splitterN246ton175n359_4 );
buf_AQFP buf_N246_splitterN246ton175n359_3_( clk_7 , buf_N246_splitterN246ton175n359_4 , 0 , buf_N246_splitterN246ton175n359_3 );
buf_AQFP buf_N246_splitterN246ton175n359_2_( clk_1 , buf_N246_splitterN246ton175n359_3 , 0 , buf_N246_splitterN246ton175n359_2 );
buf_AQFP buf_N246_splitterN246ton175n359_1_( clk_3 , buf_N246_splitterN246ton175n359_2 , 0 , buf_N246_splitterN246ton175n359_1 );
buf_AQFP buf_N260_n254_1_( clk_3 , N260 , 0 , buf_N260_n254_1 );
buf_AQFP buf_N261_splitterN261ton201n170_6_( clk_3 , N261 , 0 , buf_N261_splitterN261ton201n170_6 );
buf_AQFP buf_N261_splitterN261ton201n170_5_( clk_5 , buf_N261_splitterN261ton201n170_6 , 0 , buf_N261_splitterN261ton201n170_5 );
buf_AQFP buf_N261_splitterN261ton201n170_4_( clk_7 , buf_N261_splitterN261ton201n170_5 , 0 , buf_N261_splitterN261ton201n170_4 );
buf_AQFP buf_N261_splitterN261ton201n170_3_( clk_1 , buf_N261_splitterN261ton201n170_4 , 0 , buf_N261_splitterN261ton201n170_3 );
buf_AQFP buf_N261_splitterN261ton201n170_2_( clk_3 , buf_N261_splitterN261ton201n170_3 , 0 , buf_N261_splitterN261ton201n170_2 );
buf_AQFP buf_N261_splitterN261ton201n170_1_( clk_5 , buf_N261_splitterN261ton201n170_2 , 0 , buf_N261_splitterN261ton201n170_1 );
buf_AQFP buf_N268_splitterN268ton265n331_1_( clk_3 , N268 , 0 , buf_N268_splitterN268ton265n331_1 );
buf_AQFP buf_N55_splitterN55ton82n263_1_( clk_3 , N55 , 0 , buf_N55_splitterN55ton82n263_1 );
buf_AQFP buf_N73_n177_1_( clk_3 , N73 , 0 , buf_N73_n177_1 );
buf_AQFP buf_N74_n87_2_( clk_3 , N74 , 0 , buf_N74_n87_2 );
buf_AQFP buf_N74_n87_1_( clk_5 , buf_N74_n87_2 , 0 , buf_N74_n87_1 );
buf_AQFP buf_N80_splitterN80ton149n76_1_( clk_3 , N80 , 0 , buf_N80_splitterN80ton149n76_1 );
buf_AQFP buf_N89_n89_1_( clk_3 , N89 , 0 , buf_N89_n89_1 );
buf_AQFP buf_N90_n79_1_( clk_3 , N90 , 0 , buf_N90_n79_1 );
buf_AQFP buf_N91_splitterN91ton93n345_4_( clk_3 , N91 , 0 , buf_N91_splitterN91ton93n345_4 );
buf_AQFP buf_N91_splitterN91ton93n345_3_( clk_5 , buf_N91_splitterN91ton93n345_4 , 0 , buf_N91_splitterN91ton93n345_3 );
buf_AQFP buf_N91_splitterN91ton93n345_2_( clk_7 , buf_N91_splitterN91ton93n345_3 , 0 , buf_N91_splitterN91ton93n345_2 );
buf_AQFP buf_N91_splitterN91ton93n345_1_( clk_1 , buf_N91_splitterN91ton93n345_2 , 0 , buf_N91_splitterN91ton93n345_1 );
buf_AQFP buf_N96_splitterN96ton90n360_2_( clk_3 , N96 , 0 , buf_N96_splitterN96ton90n360_2 );
buf_AQFP buf_N96_splitterN96ton90n360_1_( clk_5 , buf_N96_splitterN96ton90n360_2 , 0 , buf_N96_splitterN96ton90n360_1 );
buf_AQFP buf_n62_N388_16_( clk_3 , n62 , 0 , buf_n62_N388_16 );
buf_AQFP buf_n62_N388_15_( clk_5 , buf_n62_N388_16 , 0 , buf_n62_N388_15 );
buf_AQFP buf_n62_N388_14_( clk_7 , buf_n62_N388_15 , 0 , buf_n62_N388_14 );
buf_AQFP buf_n62_N388_13_( clk_1 , buf_n62_N388_14 , 0 , buf_n62_N388_13 );
buf_AQFP buf_n62_N388_12_( clk_3 , buf_n62_N388_13 , 0 , buf_n62_N388_12 );
buf_AQFP buf_n62_N388_11_( clk_5 , buf_n62_N388_12 , 0 , buf_n62_N388_11 );
buf_AQFP buf_n62_N388_10_( clk_7 , buf_n62_N388_11 , 0 , buf_n62_N388_10 );
buf_AQFP buf_n62_N388_9_( clk_1 , buf_n62_N388_10 , 0 , buf_n62_N388_9 );
buf_AQFP buf_n62_N388_8_( clk_3 , buf_n62_N388_9 , 0 , buf_n62_N388_8 );
buf_AQFP buf_n62_N388_7_( clk_5 , buf_n62_N388_8 , 0 , buf_n62_N388_7 );
buf_AQFP buf_n62_N388_6_( clk_7 , buf_n62_N388_7 , 0 , buf_n62_N388_6 );
buf_AQFP buf_n62_N388_5_( clk_1 , buf_n62_N388_6 , 0 , buf_n62_N388_5 );
buf_AQFP buf_n62_N388_4_( clk_3 , buf_n62_N388_5 , 0 , buf_n62_N388_4 );
buf_AQFP buf_n62_N388_3_( clk_5 , buf_n62_N388_4 , 0 , buf_n62_N388_3 );
buf_AQFP buf_n62_N388_2_( clk_7 , buf_n62_N388_3 , 0 , buf_n62_N388_2 );
buf_AQFP buf_n62_N388_1_( clk_1 , buf_n62_N388_2 , 0 , buf_n62_N388_1 );
buf_AQFP buf_n63_splitterfromn63_1_( clk_7 , n63 , 0 , buf_n63_splitterfromn63_1 );
buf_AQFP buf_n64_N389_15_( clk_4 , n64 , 0 , buf_n64_N389_15 );
buf_AQFP buf_n64_N389_14_( clk_6 , buf_n64_N389_15 , 0 , buf_n64_N389_14 );
buf_AQFP buf_n64_N389_13_( clk_8 , buf_n64_N389_14 , 0 , buf_n64_N389_13 );
buf_AQFP buf_n64_N389_12_( clk_2 , buf_n64_N389_13 , 0 , buf_n64_N389_12 );
buf_AQFP buf_n64_N389_11_( clk_4 , buf_n64_N389_12 , 0 , buf_n64_N389_11 );
buf_AQFP buf_n64_N389_10_( clk_6 , buf_n64_N389_11 , 0 , buf_n64_N389_10 );
buf_AQFP buf_n64_N389_9_( clk_8 , buf_n64_N389_10 , 0 , buf_n64_N389_9 );
buf_AQFP buf_n64_N389_8_( clk_2 , buf_n64_N389_9 , 0 , buf_n64_N389_8 );
buf_AQFP buf_n64_N389_7_( clk_4 , buf_n64_N389_8 , 0 , buf_n64_N389_7 );
buf_AQFP buf_n64_N389_6_( clk_6 , buf_n64_N389_7 , 0 , buf_n64_N389_6 );
buf_AQFP buf_n64_N389_5_( clk_8 , buf_n64_N389_6 , 0 , buf_n64_N389_5 );
buf_AQFP buf_n64_N389_4_( clk_2 , buf_n64_N389_5 , 0 , buf_n64_N389_4 );
buf_AQFP buf_n64_N389_3_( clk_4 , buf_n64_N389_4 , 0 , buf_n64_N389_3 );
buf_AQFP buf_n64_N389_2_( clk_6 , buf_n64_N389_3 , 0 , buf_n64_N389_2 );
buf_AQFP buf_n64_N389_1_( clk_8 , buf_n64_N389_2 , 0 , buf_n64_N389_1 );
buf_AQFP buf_n65_splittern65ton72N390_13_( clk_4 , n65 , 0 , buf_n65_splittern65ton72N390_13 );
buf_AQFP buf_n65_splittern65ton72N390_12_( clk_6 , buf_n65_splittern65ton72N390_13 , 0 , buf_n65_splittern65ton72N390_12 );
buf_AQFP buf_n65_splittern65ton72N390_11_( clk_8 , buf_n65_splittern65ton72N390_12 , 0 , buf_n65_splittern65ton72N390_11 );
buf_AQFP buf_n65_splittern65ton72N390_10_( clk_2 , buf_n65_splittern65ton72N390_11 , 0 , buf_n65_splittern65ton72N390_10 );
buf_AQFP buf_n65_splittern65ton72N390_9_( clk_4 , buf_n65_splittern65ton72N390_10 , 0 , buf_n65_splittern65ton72N390_9 );
buf_AQFP buf_n65_splittern65ton72N390_8_( clk_6 , buf_n65_splittern65ton72N390_9 , 0 , buf_n65_splittern65ton72N390_8 );
buf_AQFP buf_n65_splittern65ton72N390_7_( clk_8 , buf_n65_splittern65ton72N390_8 , 0 , buf_n65_splittern65ton72N390_7 );
buf_AQFP buf_n65_splittern65ton72N390_6_( clk_2 , buf_n65_splittern65ton72N390_7 , 0 , buf_n65_splittern65ton72N390_6 );
buf_AQFP buf_n65_splittern65ton72N390_5_( clk_4 , buf_n65_splittern65ton72N390_6 , 0 , buf_n65_splittern65ton72N390_5 );
buf_AQFP buf_n65_splittern65ton72N390_4_( clk_6 , buf_n65_splittern65ton72N390_5 , 0 , buf_n65_splittern65ton72N390_4 );
buf_AQFP buf_n65_splittern65ton72N390_3_( clk_8 , buf_n65_splittern65ton72N390_4 , 0 , buf_n65_splittern65ton72N390_3 );
buf_AQFP buf_n65_splittern65ton72N390_2_( clk_2 , buf_n65_splittern65ton72N390_3 , 0 , buf_n65_splittern65ton72N390_2 );
buf_AQFP buf_n65_splittern65ton72N390_1_( clk_4 , buf_n65_splittern65ton72N390_2 , 0 , buf_n65_splittern65ton72N390_1 );
buf_AQFP buf_n66_N391_19_( clk_5 , n66 , 0 , buf_n66_N391_19 );
buf_AQFP buf_n66_N391_18_( clk_7 , buf_n66_N391_19 , 0 , buf_n66_N391_18 );
buf_AQFP buf_n66_N391_17_( clk_1 , buf_n66_N391_18 , 0 , buf_n66_N391_17 );
buf_AQFP buf_n66_N391_16_( clk_3 , buf_n66_N391_17 , 0 , buf_n66_N391_16 );
buf_AQFP buf_n66_N391_15_( clk_5 , buf_n66_N391_16 , 0 , buf_n66_N391_15 );
buf_AQFP buf_n66_N391_14_( clk_7 , buf_n66_N391_15 , 0 , buf_n66_N391_14 );
buf_AQFP buf_n66_N391_13_( clk_1 , buf_n66_N391_14 , 0 , buf_n66_N391_13 );
buf_AQFP buf_n66_N391_12_( clk_3 , buf_n66_N391_13 , 0 , buf_n66_N391_12 );
buf_AQFP buf_n66_N391_11_( clk_5 , buf_n66_N391_12 , 0 , buf_n66_N391_11 );
buf_AQFP buf_n66_N391_10_( clk_7 , buf_n66_N391_11 , 0 , buf_n66_N391_10 );
buf_AQFP buf_n66_N391_9_( clk_1 , buf_n66_N391_10 , 0 , buf_n66_N391_9 );
buf_AQFP buf_n66_N391_8_( clk_3 , buf_n66_N391_9 , 0 , buf_n66_N391_8 );
buf_AQFP buf_n66_N391_7_( clk_5 , buf_n66_N391_8 , 0 , buf_n66_N391_7 );
buf_AQFP buf_n66_N391_6_( clk_7 , buf_n66_N391_7 , 0 , buf_n66_N391_6 );
buf_AQFP buf_n66_N391_5_( clk_1 , buf_n66_N391_6 , 0 , buf_n66_N391_5 );
buf_AQFP buf_n66_N391_4_( clk_3 , buf_n66_N391_5 , 0 , buf_n66_N391_4 );
buf_AQFP buf_n66_N391_3_( clk_5 , buf_n66_N391_4 , 0 , buf_n66_N391_3 );
buf_AQFP buf_n66_N391_2_( clk_7 , buf_n66_N391_3 , 0 , buf_n66_N391_2 );
buf_AQFP buf_n66_N391_1_( clk_1 , buf_n66_N391_2 , 0 , buf_n66_N391_1 );
buf_AQFP buf_n69_N418_16_( clk_2 , n69 , 0 , buf_n69_N418_16 );
buf_AQFP buf_n69_N418_15_( clk_4 , buf_n69_N418_16 , 0 , buf_n69_N418_15 );
buf_AQFP buf_n69_N418_14_( clk_6 , buf_n69_N418_15 , 0 , buf_n69_N418_14 );
buf_AQFP buf_n69_N418_13_( clk_8 , buf_n69_N418_14 , 0 , buf_n69_N418_13 );
buf_AQFP buf_n69_N418_12_( clk_2 , buf_n69_N418_13 , 0 , buf_n69_N418_12 );
buf_AQFP buf_n69_N418_11_( clk_4 , buf_n69_N418_12 , 0 , buf_n69_N418_11 );
buf_AQFP buf_n69_N418_10_( clk_6 , buf_n69_N418_11 , 0 , buf_n69_N418_10 );
buf_AQFP buf_n69_N418_9_( clk_8 , buf_n69_N418_10 , 0 , buf_n69_N418_9 );
buf_AQFP buf_n69_N418_8_( clk_2 , buf_n69_N418_9 , 0 , buf_n69_N418_8 );
buf_AQFP buf_n69_N418_7_( clk_4 , buf_n69_N418_8 , 0 , buf_n69_N418_7 );
buf_AQFP buf_n69_N418_6_( clk_6 , buf_n69_N418_7 , 0 , buf_n69_N418_6 );
buf_AQFP buf_n69_N418_5_( clk_8 , buf_n69_N418_6 , 0 , buf_n69_N418_5 );
buf_AQFP buf_n69_N418_4_( clk_2 , buf_n69_N418_5 , 0 , buf_n69_N418_4 );
buf_AQFP buf_n69_N418_3_( clk_4 , buf_n69_N418_4 , 0 , buf_n69_N418_3 );
buf_AQFP buf_n69_N418_2_( clk_6 , buf_n69_N418_3 , 0 , buf_n69_N418_2 );
buf_AQFP buf_n69_N418_1_( clk_8 , buf_n69_N418_2 , 0 , buf_n69_N418_1 );
buf_AQFP buf_n71_splitterfromn71_14_( clk_2 , n71 , 0 , buf_n71_splitterfromn71_14 );
buf_AQFP buf_n71_splitterfromn71_13_( clk_4 , buf_n71_splitterfromn71_14 , 0 , buf_n71_splitterfromn71_13 );
buf_AQFP buf_n71_splitterfromn71_12_( clk_6 , buf_n71_splitterfromn71_13 , 0 , buf_n71_splitterfromn71_12 );
buf_AQFP buf_n71_splitterfromn71_11_( clk_8 , buf_n71_splitterfromn71_12 , 0 , buf_n71_splitterfromn71_11 );
buf_AQFP buf_n71_splitterfromn71_10_( clk_2 , buf_n71_splitterfromn71_11 , 0 , buf_n71_splitterfromn71_10 );
buf_AQFP buf_n71_splitterfromn71_9_( clk_4 , buf_n71_splitterfromn71_10 , 0 , buf_n71_splitterfromn71_9 );
buf_AQFP buf_n71_splitterfromn71_8_( clk_6 , buf_n71_splitterfromn71_9 , 0 , buf_n71_splitterfromn71_8 );
buf_AQFP buf_n71_splitterfromn71_7_( clk_8 , buf_n71_splitterfromn71_8 , 0 , buf_n71_splitterfromn71_7 );
buf_AQFP buf_n71_splitterfromn71_6_( clk_2 , buf_n71_splitterfromn71_7 , 0 , buf_n71_splitterfromn71_6 );
buf_AQFP buf_n71_splitterfromn71_5_( clk_4 , buf_n71_splitterfromn71_6 , 0 , buf_n71_splitterfromn71_5 );
buf_AQFP buf_n71_splitterfromn71_4_( clk_6 , buf_n71_splitterfromn71_5 , 0 , buf_n71_splitterfromn71_4 );
buf_AQFP buf_n71_splitterfromn71_3_( clk_8 , buf_n71_splitterfromn71_4 , 0 , buf_n71_splitterfromn71_3 );
buf_AQFP buf_n71_splitterfromn71_2_( clk_2 , buf_n71_splitterfromn71_3 , 0 , buf_n71_splitterfromn71_2 );
buf_AQFP buf_n71_splitterfromn71_1_( clk_4 , buf_n71_splitterfromn71_2 , 0 , buf_n71_splitterfromn71_1 );
buf_AQFP buf_n74_N420_15_( clk_4 , n74 , 0 , buf_n74_N420_15 );
buf_AQFP buf_n74_N420_14_( clk_6 , buf_n74_N420_15 , 0 , buf_n74_N420_14 );
buf_AQFP buf_n74_N420_13_( clk_8 , buf_n74_N420_14 , 0 , buf_n74_N420_13 );
buf_AQFP buf_n74_N420_12_( clk_2 , buf_n74_N420_13 , 0 , buf_n74_N420_12 );
buf_AQFP buf_n74_N420_11_( clk_4 , buf_n74_N420_12 , 0 , buf_n74_N420_11 );
buf_AQFP buf_n74_N420_10_( clk_6 , buf_n74_N420_11 , 0 , buf_n74_N420_10 );
buf_AQFP buf_n74_N420_9_( clk_8 , buf_n74_N420_10 , 0 , buf_n74_N420_9 );
buf_AQFP buf_n74_N420_8_( clk_2 , buf_n74_N420_9 , 0 , buf_n74_N420_8 );
buf_AQFP buf_n74_N420_7_( clk_4 , buf_n74_N420_8 , 0 , buf_n74_N420_7 );
buf_AQFP buf_n74_N420_6_( clk_6 , buf_n74_N420_7 , 0 , buf_n74_N420_6 );
buf_AQFP buf_n74_N420_5_( clk_8 , buf_n74_N420_6 , 0 , buf_n74_N420_5 );
buf_AQFP buf_n74_N420_4_( clk_2 , buf_n74_N420_5 , 0 , buf_n74_N420_4 );
buf_AQFP buf_n74_N420_3_( clk_4 , buf_n74_N420_4 , 0 , buf_n74_N420_3 );
buf_AQFP buf_n74_N420_2_( clk_6 , buf_n74_N420_3 , 0 , buf_n74_N420_2 );
buf_AQFP buf_n74_N420_1_( clk_8 , buf_n74_N420_2 , 0 , buf_n74_N420_1 );
buf_AQFP buf_n75_splitterfromn75_1_( clk_7 , n75 , 0 , buf_n75_splitterfromn75_1 );
buf_AQFP buf_n76_N421_15_( clk_4 , n76 , 0 , buf_n76_N421_15 );
buf_AQFP buf_n76_N421_14_( clk_6 , buf_n76_N421_15 , 0 , buf_n76_N421_14 );
buf_AQFP buf_n76_N421_13_( clk_8 , buf_n76_N421_14 , 0 , buf_n76_N421_13 );
buf_AQFP buf_n76_N421_12_( clk_2 , buf_n76_N421_13 , 0 , buf_n76_N421_12 );
buf_AQFP buf_n76_N421_11_( clk_4 , buf_n76_N421_12 , 0 , buf_n76_N421_11 );
buf_AQFP buf_n76_N421_10_( clk_6 , buf_n76_N421_11 , 0 , buf_n76_N421_10 );
buf_AQFP buf_n76_N421_9_( clk_8 , buf_n76_N421_10 , 0 , buf_n76_N421_9 );
buf_AQFP buf_n76_N421_8_( clk_2 , buf_n76_N421_9 , 0 , buf_n76_N421_8 );
buf_AQFP buf_n76_N421_7_( clk_4 , buf_n76_N421_8 , 0 , buf_n76_N421_7 );
buf_AQFP buf_n76_N421_6_( clk_6 , buf_n76_N421_7 , 0 , buf_n76_N421_6 );
buf_AQFP buf_n76_N421_5_( clk_8 , buf_n76_N421_6 , 0 , buf_n76_N421_5 );
buf_AQFP buf_n76_N421_4_( clk_2 , buf_n76_N421_5 , 0 , buf_n76_N421_4 );
buf_AQFP buf_n76_N421_3_( clk_4 , buf_n76_N421_4 , 0 , buf_n76_N421_3 );
buf_AQFP buf_n76_N421_2_( clk_6 , buf_n76_N421_3 , 0 , buf_n76_N421_2 );
buf_AQFP buf_n76_N421_1_( clk_8 , buf_n76_N421_2 , 0 , buf_n76_N421_1 );
buf_AQFP buf_n77_N422_15_( clk_4 , n77 , 0 , buf_n77_N422_15 );
buf_AQFP buf_n77_N422_14_( clk_6 , buf_n77_N422_15 , 0 , buf_n77_N422_14 );
buf_AQFP buf_n77_N422_13_( clk_8 , buf_n77_N422_14 , 0 , buf_n77_N422_13 );
buf_AQFP buf_n77_N422_12_( clk_2 , buf_n77_N422_13 , 0 , buf_n77_N422_12 );
buf_AQFP buf_n77_N422_11_( clk_4 , buf_n77_N422_12 , 0 , buf_n77_N422_11 );
buf_AQFP buf_n77_N422_10_( clk_6 , buf_n77_N422_11 , 0 , buf_n77_N422_10 );
buf_AQFP buf_n77_N422_9_( clk_8 , buf_n77_N422_10 , 0 , buf_n77_N422_9 );
buf_AQFP buf_n77_N422_8_( clk_2 , buf_n77_N422_9 , 0 , buf_n77_N422_8 );
buf_AQFP buf_n77_N422_7_( clk_4 , buf_n77_N422_8 , 0 , buf_n77_N422_7 );
buf_AQFP buf_n77_N422_6_( clk_6 , buf_n77_N422_7 , 0 , buf_n77_N422_6 );
buf_AQFP buf_n77_N422_5_( clk_8 , buf_n77_N422_6 , 0 , buf_n77_N422_5 );
buf_AQFP buf_n77_N422_4_( clk_2 , buf_n77_N422_5 , 0 , buf_n77_N422_4 );
buf_AQFP buf_n77_N422_3_( clk_4 , buf_n77_N422_4 , 0 , buf_n77_N422_3 );
buf_AQFP buf_n77_N422_2_( clk_6 , buf_n77_N422_3 , 0 , buf_n77_N422_2 );
buf_AQFP buf_n77_N422_1_( clk_8 , buf_n77_N422_2 , 0 , buf_n77_N422_1 );
buf_AQFP buf_n79_N423_18_( clk_6 , n79 , 0 , buf_n79_N423_18 );
buf_AQFP buf_n79_N423_17_( clk_8 , buf_n79_N423_18 , 0 , buf_n79_N423_17 );
buf_AQFP buf_n79_N423_16_( clk_2 , buf_n79_N423_17 , 0 , buf_n79_N423_16 );
buf_AQFP buf_n79_N423_15_( clk_4 , buf_n79_N423_16 , 0 , buf_n79_N423_15 );
buf_AQFP buf_n79_N423_14_( clk_6 , buf_n79_N423_15 , 0 , buf_n79_N423_14 );
buf_AQFP buf_n79_N423_13_( clk_8 , buf_n79_N423_14 , 0 , buf_n79_N423_13 );
buf_AQFP buf_n79_N423_12_( clk_2 , buf_n79_N423_13 , 0 , buf_n79_N423_12 );
buf_AQFP buf_n79_N423_11_( clk_4 , buf_n79_N423_12 , 0 , buf_n79_N423_11 );
buf_AQFP buf_n79_N423_10_( clk_6 , buf_n79_N423_11 , 0 , buf_n79_N423_10 );
buf_AQFP buf_n79_N423_9_( clk_8 , buf_n79_N423_10 , 0 , buf_n79_N423_9 );
buf_AQFP buf_n79_N423_8_( clk_2 , buf_n79_N423_9 , 0 , buf_n79_N423_8 );
buf_AQFP buf_n79_N423_7_( clk_4 , buf_n79_N423_8 , 0 , buf_n79_N423_7 );
buf_AQFP buf_n79_N423_6_( clk_6 , buf_n79_N423_7 , 0 , buf_n79_N423_6 );
buf_AQFP buf_n79_N423_5_( clk_8 , buf_n79_N423_6 , 0 , buf_n79_N423_5 );
buf_AQFP buf_n79_N423_4_( clk_2 , buf_n79_N423_5 , 0 , buf_n79_N423_4 );
buf_AQFP buf_n79_N423_3_( clk_4 , buf_n79_N423_4 , 0 , buf_n79_N423_3 );
buf_AQFP buf_n79_N423_2_( clk_6 , buf_n79_N423_3 , 0 , buf_n79_N423_2 );
buf_AQFP buf_n79_N423_1_( clk_8 , buf_n79_N423_2 , 0 , buf_n79_N423_1 );
buf_AQFP buf_n84_n85_1_( clk_7 , n84 , 0 , buf_n84_n85_1 );
buf_AQFP buf_n85_N448_16_( clk_2 , n85 , 0 , buf_n85_N448_16 );
buf_AQFP buf_n85_N448_15_( clk_4 , buf_n85_N448_16 , 0 , buf_n85_N448_15 );
buf_AQFP buf_n85_N448_14_( clk_6 , buf_n85_N448_15 , 0 , buf_n85_N448_14 );
buf_AQFP buf_n85_N448_13_( clk_8 , buf_n85_N448_14 , 0 , buf_n85_N448_13 );
buf_AQFP buf_n85_N448_12_( clk_2 , buf_n85_N448_13 , 0 , buf_n85_N448_12 );
buf_AQFP buf_n85_N448_11_( clk_4 , buf_n85_N448_12 , 0 , buf_n85_N448_11 );
buf_AQFP buf_n85_N448_10_( clk_6 , buf_n85_N448_11 , 0 , buf_n85_N448_10 );
buf_AQFP buf_n85_N448_9_( clk_8 , buf_n85_N448_10 , 0 , buf_n85_N448_9 );
buf_AQFP buf_n85_N448_8_( clk_2 , buf_n85_N448_9 , 0 , buf_n85_N448_8 );
buf_AQFP buf_n85_N448_7_( clk_4 , buf_n85_N448_8 , 0 , buf_n85_N448_7 );
buf_AQFP buf_n85_N448_6_( clk_6 , buf_n85_N448_7 , 0 , buf_n85_N448_6 );
buf_AQFP buf_n85_N448_5_( clk_8 , buf_n85_N448_6 , 0 , buf_n85_N448_5 );
buf_AQFP buf_n85_N448_4_( clk_2 , buf_n85_N448_5 , 0 , buf_n85_N448_4 );
buf_AQFP buf_n85_N448_3_( clk_4 , buf_n85_N448_4 , 0 , buf_n85_N448_3 );
buf_AQFP buf_n85_N448_2_( clk_6 , buf_n85_N448_3 , 0 , buf_n85_N448_2 );
buf_AQFP buf_n85_N448_1_( clk_8 , buf_n85_N448_2 , 0 , buf_n85_N448_1 );
buf_AQFP buf_n88_N449_16_( clk_2 , n88 , 0 , buf_n88_N449_16 );
buf_AQFP buf_n88_N449_15_( clk_4 , buf_n88_N449_16 , 0 , buf_n88_N449_15 );
buf_AQFP buf_n88_N449_14_( clk_6 , buf_n88_N449_15 , 0 , buf_n88_N449_14 );
buf_AQFP buf_n88_N449_13_( clk_8 , buf_n88_N449_14 , 0 , buf_n88_N449_13 );
buf_AQFP buf_n88_N449_12_( clk_2 , buf_n88_N449_13 , 0 , buf_n88_N449_12 );
buf_AQFP buf_n88_N449_11_( clk_4 , buf_n88_N449_12 , 0 , buf_n88_N449_11 );
buf_AQFP buf_n88_N449_10_( clk_6 , buf_n88_N449_11 , 0 , buf_n88_N449_10 );
buf_AQFP buf_n88_N449_9_( clk_8 , buf_n88_N449_10 , 0 , buf_n88_N449_9 );
buf_AQFP buf_n88_N449_8_( clk_2 , buf_n88_N449_9 , 0 , buf_n88_N449_8 );
buf_AQFP buf_n88_N449_7_( clk_4 , buf_n88_N449_8 , 0 , buf_n88_N449_7 );
buf_AQFP buf_n88_N449_6_( clk_6 , buf_n88_N449_7 , 0 , buf_n88_N449_6 );
buf_AQFP buf_n88_N449_5_( clk_8 , buf_n88_N449_6 , 0 , buf_n88_N449_5 );
buf_AQFP buf_n88_N449_4_( clk_2 , buf_n88_N449_5 , 0 , buf_n88_N449_4 );
buf_AQFP buf_n88_N449_3_( clk_4 , buf_n88_N449_4 , 0 , buf_n88_N449_3 );
buf_AQFP buf_n88_N449_2_( clk_6 , buf_n88_N449_3 , 0 , buf_n88_N449_2 );
buf_AQFP buf_n88_N449_1_( clk_8 , buf_n88_N449_2 , 0 , buf_n88_N449_1 );
buf_AQFP buf_n89_N450_18_( clk_6 , n89 , 0 , buf_n89_N450_18 );
buf_AQFP buf_n89_N450_17_( clk_8 , buf_n89_N450_18 , 0 , buf_n89_N450_17 );
buf_AQFP buf_n89_N450_16_( clk_2 , buf_n89_N450_17 , 0 , buf_n89_N450_16 );
buf_AQFP buf_n89_N450_15_( clk_4 , buf_n89_N450_16 , 0 , buf_n89_N450_15 );
buf_AQFP buf_n89_N450_14_( clk_6 , buf_n89_N450_15 , 0 , buf_n89_N450_14 );
buf_AQFP buf_n89_N450_13_( clk_8 , buf_n89_N450_14 , 0 , buf_n89_N450_13 );
buf_AQFP buf_n89_N450_12_( clk_2 , buf_n89_N450_13 , 0 , buf_n89_N450_12 );
buf_AQFP buf_n89_N450_11_( clk_4 , buf_n89_N450_12 , 0 , buf_n89_N450_11 );
buf_AQFP buf_n89_N450_10_( clk_6 , buf_n89_N450_11 , 0 , buf_n89_N450_10 );
buf_AQFP buf_n89_N450_9_( clk_8 , buf_n89_N450_10 , 0 , buf_n89_N450_9 );
buf_AQFP buf_n89_N450_8_( clk_2 , buf_n89_N450_9 , 0 , buf_n89_N450_8 );
buf_AQFP buf_n89_N450_7_( clk_4 , buf_n89_N450_8 , 0 , buf_n89_N450_7 );
buf_AQFP buf_n89_N450_6_( clk_6 , buf_n89_N450_7 , 0 , buf_n89_N450_6 );
buf_AQFP buf_n89_N450_5_( clk_8 , buf_n89_N450_6 , 0 , buf_n89_N450_5 );
buf_AQFP buf_n89_N450_4_( clk_2 , buf_n89_N450_5 , 0 , buf_n89_N450_4 );
buf_AQFP buf_n89_N450_3_( clk_4 , buf_n89_N450_4 , 0 , buf_n89_N450_3 );
buf_AQFP buf_n89_N450_2_( clk_6 , buf_n89_N450_3 , 0 , buf_n89_N450_2 );
buf_AQFP buf_n89_N450_1_( clk_8 , buf_n89_N450_2 , 0 , buf_n89_N450_1 );
buf_AQFP buf_n116_N767_10_( clk_7 , n116 , 0 , buf_n116_N767_10 );
buf_AQFP buf_n116_N767_9_( clk_1 , buf_n116_N767_10 , 0 , buf_n116_N767_9 );
buf_AQFP buf_n116_N767_8_( clk_3 , buf_n116_N767_9 , 0 , buf_n116_N767_8 );
buf_AQFP buf_n116_N767_7_( clk_5 , buf_n116_N767_8 , 0 , buf_n116_N767_7 );
buf_AQFP buf_n116_N767_6_( clk_7 , buf_n116_N767_7 , 0 , buf_n116_N767_6 );
buf_AQFP buf_n116_N767_5_( clk_1 , buf_n116_N767_6 , 0 , buf_n116_N767_5 );
buf_AQFP buf_n116_N767_4_( clk_3 , buf_n116_N767_5 , 0 , buf_n116_N767_4 );
buf_AQFP buf_n116_N767_3_( clk_5 , buf_n116_N767_4 , 0 , buf_n116_N767_3 );
buf_AQFP buf_n116_N767_2_( clk_7 , buf_n116_N767_3 , 0 , buf_n116_N767_2 );
buf_AQFP buf_n116_N767_1_( clk_1 , buf_n116_N767_2 , 0 , buf_n116_N767_1 );
buf_AQFP buf_n143_N768_12_( clk_3 , n143 , 0 , buf_n143_N768_12 );
buf_AQFP buf_n143_N768_11_( clk_5 , buf_n143_N768_12 , 0 , buf_n143_N768_11 );
buf_AQFP buf_n143_N768_10_( clk_7 , buf_n143_N768_11 , 0 , buf_n143_N768_10 );
buf_AQFP buf_n143_N768_9_( clk_1 , buf_n143_N768_10 , 0 , buf_n143_N768_9 );
buf_AQFP buf_n143_N768_8_( clk_3 , buf_n143_N768_9 , 0 , buf_n143_N768_8 );
buf_AQFP buf_n143_N768_7_( clk_5 , buf_n143_N768_8 , 0 , buf_n143_N768_7 );
buf_AQFP buf_n143_N768_6_( clk_7 , buf_n143_N768_7 , 0 , buf_n143_N768_6 );
buf_AQFP buf_n143_N768_5_( clk_1 , buf_n143_N768_6 , 0 , buf_n143_N768_5 );
buf_AQFP buf_n143_N768_4_( clk_3 , buf_n143_N768_5 , 0 , buf_n143_N768_4 );
buf_AQFP buf_n143_N768_3_( clk_5 , buf_n143_N768_4 , 0 , buf_n143_N768_3 );
buf_AQFP buf_n143_N768_2_( clk_7 , buf_n143_N768_3 , 0 , buf_n143_N768_2 );
buf_AQFP buf_n143_N768_1_( clk_1 , buf_n143_N768_2 , 0 , buf_n143_N768_1 );
buf_AQFP buf_n181_n183_1_( clk_5 , n181 , 0 , buf_n181_n183_1 );
buf_AQFP buf_n183_n184_2_( clk_8 , n183 , 0 , buf_n183_n184_2 );
buf_AQFP buf_n183_n184_1_( clk_2 , buf_n183_n184_2 , 0 , buf_n183_n184_1 );
buf_AQFP buf_n184_n185_2_( clk_5 , n184 , 0 , buf_n184_n185_2 );
buf_AQFP buf_n184_n185_1_( clk_7 , buf_n184_n185_2 , 0 , buf_n184_n185_1 );
buf_AQFP buf_n188_N850_9_( clk_8 , n188 , 0 , buf_n188_N850_9 );
buf_AQFP buf_n188_N850_8_( clk_2 , buf_n188_N850_9 , 0 , buf_n188_N850_8 );
buf_AQFP buf_n188_N850_7_( clk_4 , buf_n188_N850_8 , 0 , buf_n188_N850_7 );
buf_AQFP buf_n188_N850_6_( clk_6 , buf_n188_N850_7 , 0 , buf_n188_N850_6 );
buf_AQFP buf_n188_N850_5_( clk_8 , buf_n188_N850_6 , 0 , buf_n188_N850_5 );
buf_AQFP buf_n188_N850_4_( clk_2 , buf_n188_N850_5 , 0 , buf_n188_N850_4 );
buf_AQFP buf_n188_N850_3_( clk_4 , buf_n188_N850_4 , 0 , buf_n188_N850_3 );
buf_AQFP buf_n188_N850_2_( clk_6 , buf_n188_N850_3 , 0 , buf_n188_N850_2 );
buf_AQFP buf_n188_N850_1_( clk_8 , buf_n188_N850_2 , 0 , buf_n188_N850_1 );
buf_AQFP buf_n224_n225_2_( clk_4 , n224 , 0 , buf_n224_n225_2 );
buf_AQFP buf_n224_n225_1_( clk_6 , buf_n224_n225_2 , 0 , buf_n224_n225_1 );
buf_AQFP buf_n226_n227_1_( clk_4 , n226 , 0 , buf_n226_n227_1 );
buf_AQFP buf_n227_N863_5_( clk_8 , n227 , 0 , buf_n227_N863_5 );
buf_AQFP buf_n227_N863_4_( clk_2 , buf_n227_N863_5 , 0 , buf_n227_N863_4 );
buf_AQFP buf_n227_N863_3_( clk_4 , buf_n227_N863_4 , 0 , buf_n227_N863_3 );
buf_AQFP buf_n227_N863_2_( clk_6 , buf_n227_N863_3 , 0 , buf_n227_N863_2 );
buf_AQFP buf_n227_N863_1_( clk_8 , buf_n227_N863_2 , 0 , buf_n227_N863_1 );
buf_AQFP buf_n238_n239_1_( clk_5 , n238 , 0 , buf_n238_n239_1 );
buf_AQFP buf_n239_n240_2_( clk_8 , n239 , 0 , buf_n239_n240_2 );
buf_AQFP buf_n239_n240_1_( clk_2 , buf_n239_n240_2 , 0 , buf_n239_n240_1 );
buf_AQFP buf_n240_n241_2_( clk_5 , n240 , 0 , buf_n240_n241_2 );
buf_AQFP buf_n240_n241_1_( clk_7 , buf_n240_n241_2 , 0 , buf_n240_n241_1 );
buf_AQFP buf_n241_n242_2_( clk_3 , n241 , 0 , buf_n241_n242_2 );
buf_AQFP buf_n241_n242_1_( clk_5 , buf_n241_n242_2 , 0 , buf_n241_n242_1 );
buf_AQFP buf_n243_n244_1_( clk_3 , n243 , 0 , buf_n243_n244_1 );
buf_AQFP buf_n244_N864_6_( clk_6 , n244 , 0 , buf_n244_N864_6 );
buf_AQFP buf_n244_N864_5_( clk_8 , buf_n244_N864_6 , 0 , buf_n244_N864_5 );
buf_AQFP buf_n244_N864_4_( clk_2 , buf_n244_N864_5 , 0 , buf_n244_N864_4 );
buf_AQFP buf_n244_N864_3_( clk_4 , buf_n244_N864_4 , 0 , buf_n244_N864_3 );
buf_AQFP buf_n244_N864_2_( clk_6 , buf_n244_N864_3 , 0 , buf_n244_N864_2 );
buf_AQFP buf_n244_N864_1_( clk_8 , buf_n244_N864_2 , 0 , buf_n244_N864_1 );
buf_AQFP buf_n256_n257_2_( clk_8 , n256 , 0 , buf_n256_n257_2 );
buf_AQFP buf_n256_n257_1_( clk_2 , buf_n256_n257_2 , 0 , buf_n256_n257_1 );
buf_AQFP buf_n257_n258_2_( clk_5 , n257 , 0 , buf_n257_n258_2 );
buf_AQFP buf_n257_n258_1_( clk_7 , buf_n257_n258_2 , 0 , buf_n257_n258_1 );
buf_AQFP buf_n258_n259_1_( clk_3 , n258 , 0 , buf_n258_n259_1 );
buf_AQFP buf_n260_n261_1_( clk_8 , n260 , 0 , buf_n260_n261_1 );
buf_AQFP buf_n261_N865_8_( clk_3 , n261 , 0 , buf_n261_N865_8 );
buf_AQFP buf_n261_N865_7_( clk_5 , buf_n261_N865_8 , 0 , buf_n261_N865_7 );
buf_AQFP buf_n261_N865_6_( clk_7 , buf_n261_N865_7 , 0 , buf_n261_N865_6 );
buf_AQFP buf_n261_N865_5_( clk_1 , buf_n261_N865_6 , 0 , buf_n261_N865_5 );
buf_AQFP buf_n261_N865_4_( clk_3 , buf_n261_N865_5 , 0 , buf_n261_N865_4 );
buf_AQFP buf_n261_N865_3_( clk_5 , buf_n261_N865_4 , 0 , buf_n261_N865_3 );
buf_AQFP buf_n261_N865_2_( clk_7 , buf_n261_N865_3 , 0 , buf_n261_N865_2 );
buf_AQFP buf_n261_N865_1_( clk_1 , buf_n261_N865_2 , 0 , buf_n261_N865_1 );
buf_AQFP buf_n271_splittern271ton328n306_3_( clk_7 , n271 , 0 , buf_n271_splittern271ton328n306_3 );
buf_AQFP buf_n271_splittern271ton328n306_2_( clk_1 , buf_n271_splittern271ton328n306_3 , 0 , buf_n271_splittern271ton328n306_2 );
buf_AQFP buf_n271_splittern271ton328n306_1_( clk_3 , buf_n271_splittern271ton328n306_2 , 0 , buf_n271_splittern271ton328n306_1 );
buf_AQFP buf_n272_splitterfromn272_3_( clk_7 , n272 , 0 , buf_n272_splitterfromn272_3 );
buf_AQFP buf_n272_splitterfromn272_2_( clk_1 , buf_n272_splitterfromn272_3 , 0 , buf_n272_splitterfromn272_2 );
buf_AQFP buf_n272_splitterfromn272_1_( clk_3 , buf_n272_splitterfromn272_2 , 0 , buf_n272_splitterfromn272_1 );
buf_AQFP buf_n279_splittern279ton343n304_2_( clk_7 , n279 , 0 , buf_n279_splittern279ton343n304_2 );
buf_AQFP buf_n279_splittern279ton343n304_1_( clk_1 , buf_n279_splittern279ton343n304_2 , 0 , buf_n279_splittern279ton343n304_1 );
buf_AQFP buf_n280_splitterfromn280_3_( clk_7 , n280 , 0 , buf_n280_splitterfromn280_3 );
buf_AQFP buf_n280_splitterfromn280_2_( clk_1 , buf_n280_splitterfromn280_3 , 0 , buf_n280_splitterfromn280_2 );
buf_AQFP buf_n280_splitterfromn280_1_( clk_3 , buf_n280_splitterfromn280_2 , 0 , buf_n280_splitterfromn280_1 );
buf_AQFP buf_n287_splittern287ton358n302_1_( clk_7 , n287 , 0 , buf_n287_splittern287ton358n302_1 );
buf_AQFP buf_n288_splitterfromn288_2_( clk_7 , n288 , 0 , buf_n288_splitterfromn288_2 );
buf_AQFP buf_n288_splitterfromn288_1_( clk_1 , buf_n288_splitterfromn288_2 , 0 , buf_n288_splitterfromn288_1 );
buf_AQFP buf_n291_n292_1_( clk_2 , n291 , 0 , buf_n291_n292_1 );
buf_AQFP buf_n295_splittern295ton313n300_1_( clk_7 , n295 , 0 , buf_n295_splittern295ton313n300_1 );
buf_AQFP buf_n296_splitterfromn296_1_( clk_7 , n296 , 0 , buf_n296_splitterfromn296_1 );
buf_AQFP buf_n306_N866_1_( clk_1 , n306 , 0 , buf_n306_N866_1 );
buf_AQFP buf_n317_n318_1_( clk_1 , n317 , 0 , buf_n317_n318_1 );
buf_AQFP buf_n318_n319_4_( clk_5 , n318 , 0 , buf_n318_n319_4 );
buf_AQFP buf_n318_n319_3_( clk_7 , buf_n318_n319_4 , 0 , buf_n318_n319_3 );
buf_AQFP buf_n318_n319_2_( clk_1 , buf_n318_n319_3 , 0 , buf_n318_n319_2 );
buf_AQFP buf_n318_n319_1_( clk_3 , buf_n318_n319_2 , 0 , buf_n318_n319_1 );
buf_AQFP buf_n319_n320_1_( clk_6 , n319 , 0 , buf_n319_n320_1 );
buf_AQFP buf_n321_N874_4_( clk_3 , n321 , 0 , buf_n321_N874_4 );
buf_AQFP buf_n321_N874_3_( clk_5 , buf_n321_N874_4 , 0 , buf_n321_N874_3 );
buf_AQFP buf_n321_N874_2_( clk_7 , buf_n321_N874_3 , 0 , buf_n321_N874_2 );
buf_AQFP buf_n321_N874_1_( clk_1 , buf_n321_N874_2 , 0 , buf_n321_N874_1 );
buf_AQFP buf_n332_n333_1_( clk_2 , n332 , 0 , buf_n332_n333_1 );
buf_AQFP buf_n333_n334_5_( clk_5 , n333 , 0 , buf_n333_n334_5 );
buf_AQFP buf_n333_n334_4_( clk_7 , buf_n333_n334_5 , 0 , buf_n333_n334_4 );
buf_AQFP buf_n333_n334_3_( clk_1 , buf_n333_n334_4 , 0 , buf_n333_n334_3 );
buf_AQFP buf_n333_n334_2_( clk_3 , buf_n333_n334_3 , 0 , buf_n333_n334_2 );
buf_AQFP buf_n333_n334_1_( clk_5 , buf_n333_n334_2 , 0 , buf_n333_n334_1 );
buf_AQFP buf_n334_n335_1_( clk_1 , n334 , 0 , buf_n334_n335_1 );
buf_AQFP buf_n335_n336_2_( clk_5 , n335 , 0 , buf_n335_n336_2 );
buf_AQFP buf_n335_n336_1_( clk_7 , buf_n335_n336_2 , 0 , buf_n335_n336_1 );
buf_AQFP buf_n348_n349_5_( clk_5 , n348 , 0 , buf_n348_n349_5 );
buf_AQFP buf_n348_n349_4_( clk_7 , buf_n348_n349_5 , 0 , buf_n348_n349_4 );
buf_AQFP buf_n348_n349_3_( clk_1 , buf_n348_n349_4 , 0 , buf_n348_n349_3 );
buf_AQFP buf_n348_n349_2_( clk_3 , buf_n348_n349_3 , 0 , buf_n348_n349_2 );
buf_AQFP buf_n348_n349_1_( clk_5 , buf_n348_n349_2 , 0 , buf_n348_n349_1 );
buf_AQFP buf_n349_n350_2_( clk_8 , n349 , 0 , buf_n349_n350_2 );
buf_AQFP buf_n349_n350_1_( clk_2 , buf_n349_n350_2 , 0 , buf_n349_n350_1 );
buf_AQFP buf_n350_n351_1_( clk_5 , n350 , 0 , buf_n350_n351_1 );
buf_AQFP buf_n351_N879_1_( clk_8 , n351 , 0 , buf_n351_N879_1 );
buf_AQFP buf_n362_n363_1_( clk_2 , n362 , 0 , buf_n362_n363_1 );
buf_AQFP buf_n363_n364_4_( clk_5 , n363 , 0 , buf_n363_n364_4 );
buf_AQFP buf_n363_n364_3_( clk_7 , buf_n363_n364_4 , 0 , buf_n363_n364_3 );
buf_AQFP buf_n363_n364_2_( clk_1 , buf_n363_n364_3 , 0 , buf_n363_n364_2 );
buf_AQFP buf_n363_n364_1_( clk_3 , buf_n363_n364_2 , 0 , buf_n363_n364_1 );
buf_AQFP buf_n364_n365_1_( clk_6 , n364 , 0 , buf_n364_n365_1 );
buf_AQFP buf_n365_n366_1_( clk_2 , n365 , 0 , buf_n365_n366_1 );
buf_AQFP buf_n366_N880_3_( clk_5 , n366 , 0 , buf_n366_N880_3 );
buf_AQFP buf_n366_N880_2_( clk_7 , buf_n366_N880_3 , 0 , buf_n366_N880_2 );
buf_AQFP buf_n366_N880_1_( clk_1 , buf_n366_N880_2 , 0 , buf_n366_N880_1 );
buf_AQFP buf_splitterN1ton70n147_n147_3_( clk_4 , splitterN1ton70n147 , 0 , buf_splitterN1ton70n147_n147_3 );
buf_AQFP buf_splitterN1ton70n147_n147_2_( clk_6 , buf_splitterN1ton70n147_n147_3 , 0 , buf_splitterN1ton70n147_n147_2 );
buf_AQFP buf_splitterN1ton70n147_n147_1_( clk_8 , buf_splitterN1ton70n147_n147_2 , 0 , buf_splitterN1ton70n147_n147_1 );
buf_AQFP buf_splitterN101ton102n316_splitterN101ton281n316_3_( clk_6 , splitterN101ton102n316 , 0 , buf_splitterN101ton102n316_splitterN101ton281n316_3 );
buf_AQFP buf_splitterN101ton102n316_splitterN101ton281n316_2_( clk_8 , buf_splitterN101ton102n316_splitterN101ton281n316_3 , 0 , buf_splitterN101ton102n316_splitterN101ton281n316_2 );
buf_AQFP buf_splitterN101ton102n316_splitterN101ton281n316_1_( clk_2 , buf_splitterN101ton102n316_splitterN101ton281n316_2 , 0 , buf_splitterN101ton102n316_splitterN101ton281n316_1 );
buf_AQFP buf_splitterN106ton102n222_splitterN106ton289n222_3_( clk_5 , splitterN106ton102n222 , 0 , buf_splitterN106ton102n222_splitterN106ton289n222_3 );
buf_AQFP buf_splitterN106ton102n222_splitterN106ton289n222_2_( clk_7 , buf_splitterN106ton102n222_splitterN106ton289n222_3 , 0 , buf_splitterN106ton102n222_splitterN106ton289n222_2 );
buf_AQFP buf_splitterN106ton102n222_splitterN106ton289n222_1_( clk_1 , buf_splitterN106ton102n222_splitterN106ton289n222_2 , 0 , buf_splitterN106ton102n222_splitterN106ton289n222_1 );
buf_AQFP buf_splitterN106ton289n222_n222_1_( clk_5 , splitterN106ton289n222 , 0 , buf_splitterN106ton289n222_n222_1 );
buf_AQFP buf_splitterN111ton105n207_n207_3_( clk_6 , splitterN111ton105n207 , 0 , buf_splitterN111ton105n207_n207_3 );
buf_AQFP buf_splitterN111ton105n207_n207_2_( clk_8 , buf_splitterN111ton105n207_n207_3 , 0 , buf_splitterN111ton105n207_n207_2 );
buf_AQFP buf_splitterN111ton105n207_n207_1_( clk_2 , buf_splitterN111ton105n207_n207_2 , 0 , buf_splitterN111ton105n207_n207_1 );
buf_AQFP buf_splitterN116ton105n190_n190_3_( clk_6 , splitterN116ton105n190 , 0 , buf_splitterN116ton105n190_n190_3 );
buf_AQFP buf_splitterN116ton105n190_n190_2_( clk_8 , buf_splitterN116ton105n190_n190_3 , 0 , buf_splitterN116ton105n190_n190_2 );
buf_AQFP buf_splitterN116ton105n190_n190_1_( clk_2 , buf_splitterN116ton105n190_n190_2 , 0 , buf_splitterN116ton105n190_n190_1 );
buf_AQFP buf_splitterN121ton182n196_n196_3_( clk_5 , splitterN121ton182n196 , 0 , buf_splitterN121ton182n196_n196_3 );
buf_AQFP buf_splitterN121ton182n196_n196_2_( clk_7 , buf_splitterN121ton182n196_n196_3 , 0 , buf_splitterN121ton182n196_n196_2 );
buf_AQFP buf_splitterN121ton182n196_n196_1_( clk_1 , buf_splitterN121ton182n196_n196_2 , 0 , buf_splitterN121ton182n196_n196_1 );
buf_AQFP buf_splitterN126ton100n163_n163_1_( clk_1 , splitterN126ton100n163 , 0 , buf_splitterN126ton100n163_n163_1 );
buf_AQFP buf_splitterfromN13_n68_1_( clk_5 , splitterfromN13 , 0 , buf_splitterfromN13_n68_1 );
buf_AQFP buf_splitterfromN146_n189_1_( clk_3 , splitterfromN146 , 0 , buf_splitterfromN146_n189_1 );
buf_AQFP buf_splitterN159ton117n272_splitterN159ton330n272_4_( clk_5 , splitterN159ton117n272 , 0 , buf_splitterN159ton117n272_splitterN159ton330n272_4 );
buf_AQFP buf_splitterN159ton117n272_splitterN159ton330n272_3_( clk_7 , buf_splitterN159ton117n272_splitterN159ton330n272_4 , 0 , buf_splitterN159ton117n272_splitterN159ton330n272_3 );
buf_AQFP buf_splitterN159ton117n272_splitterN159ton330n272_2_( clk_1 , buf_splitterN159ton117n272_splitterN159ton330n272_3 , 0 , buf_splitterN159ton117n272_splitterN159ton330n272_2 );
buf_AQFP buf_splitterN159ton117n272_splitterN159ton330n272_1_( clk_3 , buf_splitterN159ton117n272_splitterN159ton330n272_2 , 0 , buf_splitterN159ton117n272_splitterN159ton330n272_1 );
buf_AQFP buf_splitterN159ton330n272_splitterN159ton271n272_3_( clk_6 , splitterN159ton330n272 , 0 , buf_splitterN159ton330n272_splitterN159ton271n272_3 );
buf_AQFP buf_splitterN159ton330n272_splitterN159ton271n272_2_( clk_8 , buf_splitterN159ton330n272_splitterN159ton271n272_3 , 0 , buf_splitterN159ton330n272_splitterN159ton271n272_2 );
buf_AQFP buf_splitterN159ton330n272_splitterN159ton271n272_1_( clk_2 , buf_splitterN159ton330n272_splitterN159ton271n272_2 , 0 , buf_splitterN159ton330n272_splitterN159ton271n272_1 );
buf_AQFP buf_splitterN165ton129n280_splitterN165ton346n280_5_( clk_5 , splitterN165ton129n280 , 0 , buf_splitterN165ton129n280_splitterN165ton346n280_5 );
buf_AQFP buf_splitterN165ton129n280_splitterN165ton346n280_4_( clk_7 , buf_splitterN165ton129n280_splitterN165ton346n280_5 , 0 , buf_splitterN165ton129n280_splitterN165ton346n280_4 );
buf_AQFP buf_splitterN165ton129n280_splitterN165ton346n280_3_( clk_1 , buf_splitterN165ton129n280_splitterN165ton346n280_4 , 0 , buf_splitterN165ton129n280_splitterN165ton346n280_3 );
buf_AQFP buf_splitterN165ton129n280_splitterN165ton346n280_2_( clk_3 , buf_splitterN165ton129n280_splitterN165ton346n280_3 , 0 , buf_splitterN165ton129n280_splitterN165ton346n280_2 );
buf_AQFP buf_splitterN165ton129n280_splitterN165ton346n280_1_( clk_5 , buf_splitterN165ton129n280_splitterN165ton346n280_2 , 0 , buf_splitterN165ton129n280_splitterN165ton346n280_1 );
buf_AQFP buf_splitterN165ton346n280_splitterN165ton279n280_2_( clk_8 , splitterN165ton346n280 , 0 , buf_splitterN165ton346n280_splitterN165ton279n280_2 );
buf_AQFP buf_splitterN165ton346n280_splitterN165ton279n280_1_( clk_2 , buf_splitterN165ton346n280_splitterN165ton279n280_2 , 0 , buf_splitterN165ton346n280_splitterN165ton279n280_1 );
buf_AQFP buf_splitterN171ton132n288_splitterN171ton361n288_4_( clk_5 , splitterN171ton132n288 , 0 , buf_splitterN171ton132n288_splitterN171ton361n288_4 );
buf_AQFP buf_splitterN171ton132n288_splitterN171ton361n288_3_( clk_7 , buf_splitterN171ton132n288_splitterN171ton361n288_4 , 0 , buf_splitterN171ton132n288_splitterN171ton361n288_3 );
buf_AQFP buf_splitterN171ton132n288_splitterN171ton361n288_2_( clk_1 , buf_splitterN171ton132n288_splitterN171ton361n288_3 , 0 , buf_splitterN171ton132n288_splitterN171ton361n288_2 );
buf_AQFP buf_splitterN171ton132n288_splitterN171ton361n288_1_( clk_3 , buf_splitterN171ton132n288_splitterN171ton361n288_2 , 0 , buf_splitterN171ton132n288_splitterN171ton361n288_1 );
buf_AQFP buf_splitterN171ton361n288_splitterN171ton287n288_2_( clk_7 , splitterN171ton361n288 , 0 , buf_splitterN171ton361n288_splitterN171ton287n288_2 );
buf_AQFP buf_splitterN171ton361n288_splitterN171ton287n288_1_( clk_1 , buf_splitterN171ton361n288_splitterN171ton287n288_2 , 0 , buf_splitterN171ton361n288_splitterN171ton287n288_1 );
buf_AQFP buf_splitterN177ton117n296_splitterN177ton315n296_3_( clk_5 , splitterN177ton117n296 , 0 , buf_splitterN177ton117n296_splitterN177ton315n296_3 );
buf_AQFP buf_splitterN177ton117n296_splitterN177ton315n296_2_( clk_7 , buf_splitterN177ton117n296_splitterN177ton315n296_3 , 0 , buf_splitterN177ton117n296_splitterN177ton315n296_2 );
buf_AQFP buf_splitterN177ton117n296_splitterN177ton315n296_1_( clk_1 , buf_splitterN177ton117n296_splitterN177ton315n296_2 , 0 , buf_splitterN177ton117n296_splitterN177ton315n296_1 );
buf_AQFP buf_splitterN177ton315n296_splitterN177ton295n296_3_( clk_5 , splitterN177ton315n296 , 0 , buf_splitterN177ton315n296_splitterN177ton295n296_3 );
buf_AQFP buf_splitterN177ton315n296_splitterN177ton295n296_2_( clk_7 , buf_splitterN177ton315n296_splitterN177ton295n296_3 , 0 , buf_splitterN177ton315n296_splitterN177ton295n296_2 );
buf_AQFP buf_splitterN177ton315n296_splitterN177ton295n296_1_( clk_1 , buf_splitterN177ton315n296_splitterN177ton295n296_2 , 0 , buf_splitterN177ton315n296_splitterN177ton295n296_1 );
buf_AQFP buf_splitterN183ton132n212_splitterN183ton221n212_4_( clk_5 , splitterN183ton132n212 , 0 , buf_splitterN183ton132n212_splitterN183ton221n212_4 );
buf_AQFP buf_splitterN183ton132n212_splitterN183ton221n212_3_( clk_7 , buf_splitterN183ton132n212_splitterN183ton221n212_4 , 0 , buf_splitterN183ton132n212_splitterN183ton221n212_3 );
buf_AQFP buf_splitterN183ton132n212_splitterN183ton221n212_2_( clk_1 , buf_splitterN183ton132n212_splitterN183ton221n212_3 , 0 , buf_splitterN183ton132n212_splitterN183ton221n212_2 );
buf_AQFP buf_splitterN183ton132n212_splitterN183ton221n212_1_( clk_3 , buf_splitterN183ton132n212_splitterN183ton221n212_2 , 0 , buf_splitterN183ton132n212_splitterN183ton221n212_1 );
buf_AQFP buf_splitterN183ton221n212_splitterN183ton211n212_2_( clk_7 , splitterN183ton221n212 , 0 , buf_splitterN183ton221n212_splitterN183ton211n212_2 );
buf_AQFP buf_splitterN183ton221n212_splitterN183ton211n212_1_( clk_1 , buf_splitterN183ton221n212_splitterN183ton211n212_2 , 0 , buf_splitterN183ton221n212_splitterN183ton211n212_1 );
buf_AQFP buf_splitterN189ton123n194_splitterN189ton236n194_2_( clk_5 , splitterN189ton123n194 , 0 , buf_splitterN189ton123n194_splitterN189ton236n194_2 );
buf_AQFP buf_splitterN189ton123n194_splitterN189ton236n194_1_( clk_7 , buf_splitterN189ton123n194_splitterN189ton236n194_2 , 0 , buf_splitterN189ton123n194_splitterN189ton236n194_1 );
buf_AQFP buf_splitterN189ton236n194_splitterN189ton193n194_3_( clk_3 , splitterN189ton236n194 , 0 , buf_splitterN189ton236n194_splitterN189ton193n194_3 );
buf_AQFP buf_splitterN189ton236n194_splitterN189ton193n194_2_( clk_5 , buf_splitterN189ton236n194_splitterN189ton193n194_3 , 0 , buf_splitterN189ton236n194_splitterN189ton193n194_2 );
buf_AQFP buf_splitterN189ton236n194_splitterN189ton193n194_1_( clk_7 , buf_splitterN189ton236n194_splitterN189ton193n194_2 , 0 , buf_splitterN189ton236n194_splitterN189ton193n194_1 );
buf_AQFP buf_splitterN195ton123n200_splitterN195ton253n200_2_( clk_5 , splitterN195ton123n200 , 0 , buf_splitterN195ton123n200_splitterN195ton253n200_2 );
buf_AQFP buf_splitterN195ton123n200_splitterN195ton253n200_1_( clk_7 , buf_splitterN195ton123n200_splitterN195ton253n200_2 , 0 , buf_splitterN195ton123n200_splitterN195ton253n200_1 );
buf_AQFP buf_splitterN195ton253n200_splitterN195ton199n200_2_( clk_3 , splitterN195ton253n200 , 0 , buf_splitterN195ton253n200_splitterN195ton199n200_2 );
buf_AQFP buf_splitterN195ton253n200_splitterN195ton199n200_1_( clk_5 , buf_splitterN195ton253n200_splitterN195ton199n200_2 , 0 , buf_splitterN195ton253n200_splitterN195ton199n200_1 );
buf_AQFP buf_splitterN201ton129n167_splitterN201ton180n167_2_( clk_5 , splitterN201ton129n167 , 0 , buf_splitterN201ton129n167_splitterN201ton180n167_2 );
buf_AQFP buf_splitterN201ton129n167_splitterN201ton180n167_1_( clk_7 , buf_splitterN201ton129n167_splitterN201ton180n167_2 , 0 , buf_splitterN201ton129n167_splitterN201ton180n167_1 );
buf_AQFP buf_splitterN201ton180n167_splitterN201ton166n167_2_( clk_2 , splitterN201ton180n167 , 0 , buf_splitterN201ton180n167_splitterN201ton166n167_2 );
buf_AQFP buf_splitterN201ton180n167_splitterN201ton166n167_1_( clk_4 , buf_splitterN201ton180n167_splitterN201ton166n167_2 , 0 , buf_splitterN201ton180n167_splitterN201ton166n167_1 );
buf_AQFP buf_splitterN210ton182n345_splitterN210ton316n345_3_( clk_5 , splitterN210ton182n345 , 0 , buf_splitterN210ton182n345_splitterN210ton316n345_3 );
buf_AQFP buf_splitterN210ton182n345_splitterN210ton316n345_2_( clk_7 , buf_splitterN210ton182n345_splitterN210ton316n345_3 , 0 , buf_splitterN210ton182n345_splitterN210ton316n345_2 );
buf_AQFP buf_splitterN210ton182n345_splitterN210ton316n345_1_( clk_1 , buf_splitterN210ton182n345_splitterN210ton316n345_2 , 0 , buf_splitterN210ton182n345_splitterN210ton316n345_1 );
buf_AQFP buf_splitterN219ton171n325_splitterN219ton249n325_1_( clk_4 , splitterN219ton171n325 , 0 , buf_splitterN219ton171n325_splitterN219ton249n325_1 );
buf_AQFP buf_splitterN219ton249n325_splitterN219ton232n325_1_( clk_7 , splitterN219ton249n325 , 0 , buf_splitterN219ton249n325_splitterN219ton232n325_1 );
buf_AQFP buf_splitterN219ton232n325_splitterN219ton217n325_1_( clk_2 , splitterN219ton232n325 , 0 , buf_splitterN219ton232n325_splitterN219ton217n325_1 );
buf_AQFP buf_splitterN219ton217n325_splitterN219ton355n325_1_( clk_5 , splitterN219ton217n325 , 0 , buf_splitterN219ton217n325_splitterN219ton355n325_1 );
buf_AQFP buf_splitterN219ton355n325_splitterN219ton340n325_1_( clk_1 , splitterN219ton355n325 , 0 , buf_splitterN219ton355n325_splitterN219ton340n325_1 );
buf_AQFP buf_splitterN219ton340n325_n325_2_( clk_4 , splitterN219ton340n325 , 0 , buf_splitterN219ton340n325_n325_2 );
buf_AQFP buf_splitterN219ton340n325_n325_1_( clk_6 , buf_splitterN219ton340n325_n325_2 , 0 , buf_splitterN219ton340n325_n325_1 );
buf_AQFP buf_splitterN228ton250n342_splitterN228ton233n342_1_( clk_5 , splitterN228ton250n342 , 0 , buf_splitterN228ton250n342_splitterN228ton233n342_1 );
buf_AQFP buf_splitterN228ton218n342_splitterN228ton309n342_1_( clk_2 , splitterN228ton218n342 , 0 , buf_splitterN228ton218n342_splitterN228ton309n342_1 );
buf_AQFP buf_splitterN237ton174n328_splitterN237ton251n328_1_( clk_1 , splitterN237ton174n328 , 0 , buf_splitterN237ton174n328_splitterN237ton251n328_1 );
buf_AQFP buf_splitterN268ton265n331_splitterN268ton152n331_1_( clk_7 , splitterN268ton265n331 , 0 , buf_splitterN268ton265n331_splitterN268ton152n331_1 );
buf_AQFP buf_splitterN268ton152n331_n331_2_( clk_3 , splitterN268ton152n331 , 0 , buf_splitterN268ton152n331_n331_2 );
buf_AQFP buf_splitterN268ton152n331_n331_1_( clk_5 , buf_splitterN268ton152n331_n331_2 , 0 , buf_splitterN268ton152n331_n331_1 );
buf_AQFP buf_splitterN51ton81n275_n275_2_( clk_6 , splitterN51ton81n275 , 0 , buf_splitterN51ton81n275_n275_2 );
buf_AQFP buf_splitterN51ton81n275_n275_1_( clk_8 , buf_splitterN51ton81n275_n275_2 , 0 , buf_splitterN51ton81n275_n275_1 );
buf_AQFP buf_splitterN55ton82n263_splitterN55ton151n263_1_( clk_6 , splitterN55ton82n263 , 0 , buf_splitterN55ton82n263_splitterN55ton151n263_1 );
buf_AQFP buf_splitterfromN8_n267_2_( clk_5 , splitterfromN8 , 0 , buf_splitterfromN8_n267_2 );
buf_AQFP buf_splitterfromN8_n267_1_( clk_7 , buf_splitterfromN8_n267_2 , 0 , buf_splitterfromN8_n267_1 );
buf_AQFP buf_splitterN80ton149n76_splitterN80ton64n76_1_( clk_7 , splitterN80ton149n76 , 0 , buf_splitterN80ton149n76_splitterN80ton64n76_1 );
buf_AQFP buf_splitterN96ton90n360_splitterN96ton273n360_2_( clk_8 , splitterN96ton90n360 , 0 , buf_splitterN96ton90n360_splitterN96ton273n360_2 );
buf_AQFP buf_splitterN96ton90n360_splitterN96ton273n360_1_( clk_2 , buf_splitterN96ton90n360_splitterN96ton273n360_2 , 0 , buf_splitterN96ton90n360_splitterN96ton273n360_1 );
buf_AQFP buf_splitterN96ton273n360_n360_1_( clk_5 , splitterN96ton273n360 , 0 , buf_splitterN96ton273n360_n360_1 );
buf_AQFP buf_splitterfromn61_n62_1_( clk_7 , splitterfromn61 , 0 , buf_splitterfromn61_n62_1 );
buf_AQFP buf_splittern65ton72N390_N390_1_( clk_8 , splittern65ton72N390 , 0 , buf_splittern65ton72N390_N390_1 );
buf_AQFP buf_splittern67ton160n69_n69_1_( clk_7 , splittern67ton160n69 , 0 , buf_splittern67ton160n69_n69_1 );
buf_AQFP buf_splitterfromn70_n71_1_( clk_6 , splitterfromn70 , 0 , buf_splitterfromn70_n71_1 );
buf_AQFP buf_splitterfromn73_n74_1_( clk_8 , splitterfromn73 , 0 , buf_splitterfromn73_n74_1 );
buf_AQFP buf_splittern81ton145N447_N447_17_( clk_8 , splittern81ton145N447 , 0 , buf_splittern81ton145N447_N447_17 );
buf_AQFP buf_splittern81ton145N447_N447_16_( clk_2 , buf_splittern81ton145N447_N447_17 , 0 , buf_splittern81ton145N447_N447_16 );
buf_AQFP buf_splittern81ton145N447_N447_15_( clk_4 , buf_splittern81ton145N447_N447_16 , 0 , buf_splittern81ton145N447_N447_15 );
buf_AQFP buf_splittern81ton145N447_N447_14_( clk_6 , buf_splittern81ton145N447_N447_15 , 0 , buf_splittern81ton145N447_N447_14 );
buf_AQFP buf_splittern81ton145N447_N447_13_( clk_8 , buf_splittern81ton145N447_N447_14 , 0 , buf_splittern81ton145N447_N447_13 );
buf_AQFP buf_splittern81ton145N447_N447_12_( clk_2 , buf_splittern81ton145N447_N447_13 , 0 , buf_splittern81ton145N447_N447_12 );
buf_AQFP buf_splittern81ton145N447_N447_11_( clk_4 , buf_splittern81ton145N447_N447_12 , 0 , buf_splittern81ton145N447_N447_11 );
buf_AQFP buf_splittern81ton145N447_N447_10_( clk_6 , buf_splittern81ton145N447_N447_11 , 0 , buf_splittern81ton145N447_N447_10 );
buf_AQFP buf_splittern81ton145N447_N447_9_( clk_8 , buf_splittern81ton145N447_N447_10 , 0 , buf_splittern81ton145N447_N447_9 );
buf_AQFP buf_splittern81ton145N447_N447_8_( clk_2 , buf_splittern81ton145N447_N447_9 , 0 , buf_splittern81ton145N447_N447_8 );
buf_AQFP buf_splittern81ton145N447_N447_7_( clk_4 , buf_splittern81ton145N447_N447_8 , 0 , buf_splittern81ton145N447_N447_7 );
buf_AQFP buf_splittern81ton145N447_N447_6_( clk_6 , buf_splittern81ton145N447_N447_7 , 0 , buf_splittern81ton145N447_N447_6 );
buf_AQFP buf_splittern81ton145N447_N447_5_( clk_8 , buf_splittern81ton145N447_N447_6 , 0 , buf_splittern81ton145N447_N447_5 );
buf_AQFP buf_splittern81ton145N447_N447_4_( clk_2 , buf_splittern81ton145N447_N447_5 , 0 , buf_splittern81ton145N447_N447_4 );
buf_AQFP buf_splittern81ton145N447_N447_3_( clk_4 , buf_splittern81ton145N447_N447_4 , 0 , buf_splittern81ton145N447_N447_3 );
buf_AQFP buf_splittern81ton145N447_N447_2_( clk_6 , buf_splittern81ton145N447_N447_3 , 0 , buf_splittern81ton145N447_N447_2 );
buf_AQFP buf_splittern81ton145N447_N447_1_( clk_8 , buf_splittern81ton145N447_N447_2 , 0 , buf_splittern81ton145N447_N447_1 );
buf_AQFP buf_splittern152ton164n210_n210_1_( clk_5 , splittern152ton164n210 , 0 , buf_splittern152ton164n210_n210_1 );
buf_AQFP buf_splittern193ton228n206_n206_1_( clk_7 , splittern193ton228n206 , 0 , buf_splittern193ton228n206_n206_1 );
buf_AQFP buf_splittern199ton245n204_n204_1_( clk_4 , splittern199ton245n204 , 0 , buf_splittern199ton245n204_n204_1 );
buf_AQFP buf_splittern211ton213n298_n298_2_( clk_8 , splittern211ton213n298 , 0 , buf_splittern211ton213n298_n298_2 );
buf_AQFP buf_splittern211ton213n298_n298_1_( clk_2 , buf_splittern211ton213n298_n298_2 , 0 , buf_splittern211ton213n298_n298_1 );
buf_AQFP buf_splitterfromn212_n297_1_( clk_8 , splitterfromn212 , 0 , buf_splitterfromn212_n297_1 );
buf_AQFP buf_splittern271ton328n306_n306_4_( clk_7 , splittern271ton328n306 , 0 , buf_splittern271ton328n306_n306_4 );
buf_AQFP buf_splittern271ton328n306_n306_3_( clk_1 , buf_splittern271ton328n306_n306_4 , 0 , buf_splittern271ton328n306_n306_3 );
buf_AQFP buf_splittern271ton328n306_n306_2_( clk_3 , buf_splittern271ton328n306_n306_3 , 0 , buf_splittern271ton328n306_n306_2 );
buf_AQFP buf_splittern271ton328n306_n306_1_( clk_5 , buf_splittern271ton328n306_n306_2 , 0 , buf_splittern271ton328n306_n306_1 );
buf_AQFP buf_splitterfromn272_n305_4_( clk_7 , splitterfromn272 , 0 , buf_splitterfromn272_n305_4 );
buf_AQFP buf_splitterfromn272_n305_3_( clk_1 , buf_splitterfromn272_n305_4 , 0 , buf_splitterfromn272_n305_3 );
buf_AQFP buf_splitterfromn272_n305_2_( clk_3 , buf_splitterfromn272_n305_3 , 0 , buf_splitterfromn272_n305_2 );
buf_AQFP buf_splitterfromn272_n305_1_( clk_5 , buf_splitterfromn272_n305_2 , 0 , buf_splitterfromn272_n305_1 );
buf_AQFP buf_splittern279ton337n304_n304_3_( clk_7 , splittern279ton337n304 , 0 , buf_splittern279ton337n304_n304_3 );
buf_AQFP buf_splittern279ton337n304_n304_2_( clk_1 , buf_splittern279ton337n304_n304_3 , 0 , buf_splittern279ton337n304_n304_2 );
buf_AQFP buf_splittern279ton337n304_n304_1_( clk_3 , buf_splittern279ton337n304_n304_2 , 0 , buf_splittern279ton337n304_n304_1 );
buf_AQFP buf_splitterfromn280_n303_2_( clk_7 , splitterfromn280 , 0 , buf_splitterfromn280_n303_2 );
buf_AQFP buf_splitterfromn280_n303_1_( clk_1 , buf_splitterfromn280_n303_2 , 0 , buf_splitterfromn280_n303_1 );
buf_AQFP buf_splittern287ton352n302_n302_2_( clk_5 , splittern287ton352n302 , 0 , buf_splittern287ton352n302_n302_2 );
buf_AQFP buf_splittern287ton352n302_n302_1_( clk_7 , buf_splittern287ton352n302_n302_2 , 0 , buf_splittern287ton352n302_n302_1 );
buf_AQFP buf_splitterfromn288_n301_2_( clk_4 , splitterfromn288 , 0 , buf_splitterfromn288_n301_2 );
buf_AQFP buf_splitterfromn288_n301_1_( clk_6 , buf_splitterfromn288_n301_2 , 0 , buf_splitterfromn288_n301_1 );
buf_AQFP buf_splittern295ton313n300_n300_2_( clk_2 , splittern295ton313n300 , 0 , buf_splittern295ton313n300_n300_2 );
buf_AQFP buf_splittern295ton313n300_n300_1_( clk_4 , buf_splittern295ton313n300_n300_2 , 0 , buf_splittern295ton313n300_n300_1 );
buf_AQFP buf_splitterfromn296_n299_2_( clk_2 , splitterfromn296 , 0 , buf_splitterfromn296_n299_2 );
buf_AQFP buf_splitterfromn296_n299_1_( clk_4 , buf_splitterfromn296_n299_2 , 0 , buf_splitterfromn296_n299_1 );
buf_AQFP buf_splitterfromn307_n310_1_( clk_6 , splitterfromn307 , 0 , buf_splitterfromn307_n310_1 );
buf_AQFP buf_splittern322ton327n324_splittern322ton323n324_1_( clk_3 , splittern322ton327n324 , 0 , buf_splittern322ton327n324_splittern322ton323n324_1 );
splitter_AQFP splitterN1ton70n147_( clk_2 , N1 , 0 , splitterN1ton70n147 );
splitter_AQFP splitterN101ton102n316_( clk_4 , buf_N101_splitterN101ton102n316_1 , 0 , splitterN101ton102n316 );
splitter_AQFP splitterN101ton281n316_( clk_3 , buf_splitterN101ton102n316_splitterN101ton281n316_1 , 0 , splitterN101ton281n316 );
splitter_AQFP splitterN106ton102n222_( clk_3 , N106 , 0 , splitterN106ton102n222 );
splitter_AQFP splitterN106ton289n222_( clk_3 , buf_splitterN106ton102n222_splitterN106ton289n222_1 , 0 , splitterN106ton289n222 );
splitter_AQFP splitterN111ton105n207_( clk_4 , buf_N111_splitterN111ton105n207_1 , 0 , splitterN111ton105n207 );
splitter_AQFP splitterN116ton105n190_( clk_4 , buf_N116_splitterN116ton105n190_1 , 0 , splitterN116ton105n190 );
splitter_AQFP splitterN121ton182n196_( clk_3 , N121 , 0 , splitterN121ton182n196 );
splitter_AQFP splitterN126ton100n163_( clk_7 , buf_N126_splitterN126ton100n163_1 , 0 , splitterN126ton100n163 );
splitter_AQFP splitterfromN13_( clk_3 , N13 , 0 , splitterfromN13 );
splitter_AQFP splitterN130ton90n121_( clk_5 , buf_N130_splitterN130ton90n121_1 , 0 , splitterN130ton90n121 );
splitter_AQFP splitterN130ton120n121_( clk_7 , splitterN130ton90n121 , 0 , splitterN130ton120n121 );
splitter_AQFP splitterfromN135_( clk_2 , N135 , 0 , splitterfromN135 );
splitter_AQFP splitterN138ton291n283_( clk_7 , buf_N138_splitterN138ton291n283_1 , 0 , splitterN138ton291n283 );
splitter_AQFP splitterfromN143_( clk_2 , buf_N143_splitterfromN143_1 , 0 , splitterfromN143 );
splitter_AQFP splitterfromN146_( clk_1 , buf_N146_splitterfromN146_1 , 0 , splitterfromN146 );
splitter_AQFP splitterfromN149_( clk_2 , buf_N149_splitterfromN149_1 , 0 , splitterfromN149 );
splitter_AQFP splitterfromN153_( clk_2 , buf_N153_splitterfromN153_1 , 0 , splitterfromN153 );
splitter_AQFP splitterN159ton117n272_( clk_3 , N159 , 0 , splitterN159ton117n272 );
splitter_AQFP splitterN159ton330n272_( clk_4 , buf_splitterN159ton117n272_splitterN159ton330n272_1 , 0 , splitterN159ton330n272 );
splitter_AQFP splitterN159ton271n272_( clk_3 , buf_splitterN159ton330n272_splitterN159ton271n272_1 , 0 , splitterN159ton271n272 );
splitter_AQFP splitterN165ton129n280_( clk_3 , N165 , 0 , splitterN165ton129n280 );
splitter_AQFP splitterN165ton346n280_( clk_6 , buf_splitterN165ton129n280_splitterN165ton346n280_1 , 0 , splitterN165ton346n280 );
splitter_AQFP splitterN165ton279n280_( clk_3 , buf_splitterN165ton346n280_splitterN165ton279n280_1 , 0 , splitterN165ton279n280 );
splitter_AQFP splitterN17ton153n283_( clk_3 , N17 , 0 , splitterN17ton153n283 );
splitter_AQFP splitterN17ton68n283_( clk_5 , splitterN17ton153n283 , 0 , splitterN17ton68n283 );
splitter_AQFP splitterN17ton146n283_( clk_7 , splitterN17ton68n283 , 0 , splitterN17ton146n283 );
splitter_AQFP splitterN171ton132n288_( clk_3 , N171 , 0 , splitterN171ton132n288 );
splitter_AQFP splitterN171ton361n288_( clk_5 , buf_splitterN171ton132n288_splitterN171ton361n288_1 , 0 , splitterN171ton361n288 );
splitter_AQFP splitterN171ton287n288_( clk_3 , buf_splitterN171ton361n288_splitterN171ton287n288_1 , 0 , splitterN171ton287n288 );
splitter_AQFP splitterN177ton117n296_( clk_3 , N177 , 0 , splitterN177ton117n296 );
splitter_AQFP splitterN177ton315n296_( clk_3 , buf_splitterN177ton117n296_splitterN177ton315n296_1 , 0 , splitterN177ton315n296 );
splitter_AQFP splitterN177ton295n296_( clk_3 , buf_splitterN177ton315n296_splitterN177ton295n296_1 , 0 , splitterN177ton295n296 );
splitter_AQFP splitterN183ton132n212_( clk_3 , N183 , 0 , splitterN183ton132n212 );
splitter_AQFP splitterN183ton221n212_( clk_5 , buf_splitterN183ton132n212_splitterN183ton221n212_1 , 0 , splitterN183ton221n212 );
splitter_AQFP splitterN183ton211n212_( clk_2 , buf_splitterN183ton221n212_splitterN183ton211n212_1 , 0 , splitterN183ton211n212 );
splitter_AQFP splitterN189ton123n194_( clk_3 , N189 , 0 , splitterN189ton123n194 );
splitter_AQFP splitterN189ton236n194_( clk_1 , buf_splitterN189ton123n194_splitterN189ton236n194_1 , 0 , splitterN189ton236n194 );
splitter_AQFP splitterN189ton193n194_( clk_1 , buf_splitterN189ton236n194_splitterN189ton193n194_1 , 0 , splitterN189ton193n194 );
splitter_AQFP splitterN195ton123n200_( clk_3 , N195 , 0 , splitterN195ton123n200 );
splitter_AQFP splitterN195ton253n200_( clk_1 , buf_splitterN195ton123n200_splitterN195ton253n200_1 , 0 , splitterN195ton253n200 );
splitter_AQFP splitterN195ton199n200_( clk_6 , buf_splitterN195ton253n200_splitterN195ton199n200_1 , 0 , splitterN195ton199n200 );
splitter_AQFP splitterN201ton129n167_( clk_3 , N201 , 0 , splitterN201ton129n167 );
splitter_AQFP splitterN201ton180n167_( clk_8 , buf_splitterN201ton129n167_splitterN201ton180n167_1 , 0 , splitterN201ton180n167 );
splitter_AQFP splitterN201ton166n167_( clk_5 , buf_splitterN201ton180n167_splitterN201ton166n167_1 , 0 , splitterN201ton166n167 );
splitter_AQFP splitterfromN207_( clk_5 , buf_N207_splitterfromN207_1 , 0 , splitterfromN207 );
splitter_AQFP splitterN210ton182n345_( clk_3 , N210 , 0 , splitterN210ton182n345 );
splitter_AQFP splitterN210ton316n345_( clk_3 , buf_splitterN210ton182n345_splitterN210ton316n345_1 , 0 , splitterN210ton316n345 );
splitter_AQFP splitterN210ton222n345_( clk_5 , splitterN210ton316n345 , 0 , splitterN210ton222n345 );
splitter_AQFP splitterN219ton171n325_( clk_2 , buf_N219_splitterN219ton171n325_1 , 0 , splitterN219ton171n325 );
splitter_AQFP splitterN219ton249n325_( clk_5 , buf_splitterN219ton171n325_splitterN219ton249n325_1 , 0 , splitterN219ton249n325 );
splitter_AQFP splitterN219ton232n325_( clk_8 , buf_splitterN219ton249n325_splitterN219ton232n325_1 , 0 , splitterN219ton232n325 );
splitter_AQFP splitterN219ton217n325_( clk_3 , buf_splitterN219ton232n325_splitterN219ton217n325_1 , 0 , splitterN219ton217n325 );
splitter_AQFP splitterN219ton355n325_( clk_7 , buf_splitterN219ton217n325_splitterN219ton355n325_1 , 0 , splitterN219ton355n325 );
splitter_AQFP splitterN219ton340n325_( clk_2 , buf_splitterN219ton355n325_splitterN219ton340n325_1 , 0 , splitterN219ton340n325 );
splitter_AQFP splitterN228ton173n342_( clk_1 , buf_N228_splitterN228ton173n342_1 , 0 , splitterN228ton173n342 );
splitter_AQFP splitterN228ton250n342_( clk_3 , splitterN228ton173n342 , 0 , splitterN228ton250n342 );
splitter_AQFP splitterN228ton233n342_( clk_6 , buf_splitterN228ton250n342_splitterN228ton233n342_1 , 0 , splitterN228ton233n342 );
splitter_AQFP splitterN228ton218n342_( clk_8 , splitterN228ton233n342 , 0 , splitterN228ton218n342 );
splitter_AQFP splitterN228ton309n342_( clk_4 , buf_splitterN228ton218n342_splitterN228ton309n342_1 , 0 , splitterN228ton309n342 );
splitter_AQFP splitterN228ton357n342_( clk_6 , splitterN228ton309n342 , 0 , splitterN228ton357n342 );
splitter_AQFP splitterN228ton327n342_( clk_8 , splitterN228ton357n342 , 0 , splitterN228ton327n342 );
splitter_AQFP splitterN237ton174n328_( clk_7 , buf_N237_splitterN237ton174n328_1 , 0 , splitterN237ton174n328 );
splitter_AQFP splitterN237ton251n328_( clk_2 , buf_splitterN237ton174n328_splitterN237ton251n328_1 , 0 , splitterN237ton251n328 );
splitter_AQFP splitterN237ton234n328_( clk_4 , splitterN237ton251n328 , 0 , splitterN237ton234n328 );
splitter_AQFP splitterN237ton219n328_( clk_6 , splitterN237ton234n328 , 0 , splitterN237ton219n328 );
splitter_AQFP splitterN237ton313n328_( clk_8 , splitterN237ton219n328 , 0 , splitterN237ton313n328 );
splitter_AQFP splitterN237ton358n328_( clk_2 , splitterN237ton313n328 , 0 , splitterN237ton358n328 );
splitter_AQFP splitterN237ton343n328_( clk_4 , splitterN237ton358n328 , 0 , splitterN237ton343n328 );
splitter_AQFP splitterN246ton175n359_( clk_5 , buf_N246_splitterN246ton175n359_1 , 0 , splitterN246ton175n359 );
splitter_AQFP splitterN246ton235n359_( clk_7 , splitterN246ton175n359 , 0 , splitterN246ton235n359 );
splitter_AQFP splitterN246ton314n359_( clk_8 , splitterN246ton235n359 , 0 , splitterN246ton314n359 );
splitter_AQFP splitterN255ton181n254_( clk_2 , N255 , 0 , splitterN255ton181n254 );
splitter_AQFP splitterN261ton201n170_( clk_7 , buf_N261_splitterN261ton201n170_1 , 0 , splitterN261ton201n170 );
splitter_AQFP splitterN261ton169n170_( clk_1 , splitterN261ton201n170 , 0 , splitterN261ton169n170 );
splitter_AQFP splitterN268ton265n331_( clk_5 , buf_N268_splitterN268ton265n331_1 , 0 , splitterN268ton265n331 );
splitter_AQFP splitterN268ton152n331_( clk_1 , buf_splitterN268ton265n331_splitterN268ton152n331_1 , 0 , splitterN268ton152n331 );
splitter_AQFP splitterN29ton61n84_( clk_3 , N29 , 0 , splitterN29ton61n84 );
splitter_AQFP splitterfromN36_( clk_3 , N36 , 0 , splitterfromN36 );
splitter_AQFP splitterN42ton176n77_( clk_2 , N42 , 0 , splitterN42ton176n77 );
splitter_AQFP splitterN42ton153n77_( clk_4 , splitterN42ton176n77 , 0 , splitterN42ton153n77 );
splitter_AQFP splitterN42ton158n77_( clk_6 , splitterN42ton153n77 , 0 , splitterN42ton158n77 );
splitter_AQFP splitterN42ton62n77_( clk_8 , splitterN42ton158n77 , 0 , splitterN42ton62n77 );
splitter_AQFP splitterN51ton159n275_( clk_3 , N51 , 0 , splitterN51ton159n275 );
splitter_AQFP splitterN51ton81n275_( clk_4 , splitterN51ton159n275 , 0 , splitterN51ton81n275 );
splitter_AQFP splitterN55ton82n263_( clk_4 , buf_N55_splitterN55ton82n263_1 , 0 , splitterN55ton82n263 );
splitter_AQFP splitterN55ton151n263_( clk_7 , buf_splitterN55ton82n263_splitterN55ton151n263_1 , 0 , splitterN55ton151n263 );
splitter_AQFP splitterN59ton144n75_( clk_2 , N59 , 0 , splitterN59ton144n75 );
splitter_AQFP splitterN59ton73n75_( clk_3 , splitterN59ton144n75 , 0 , splitterN59ton73n75 );
splitter_AQFP splitterfromN68_( clk_3 , N68 , 0 , splitterfromN68 );
splitter_AQFP splitterfromN75_( clk_3 , N75 , 0 , splitterfromN75 );
splitter_AQFP splitterfromN8_( clk_3 , N8 , 0 , splitterfromN8 );
splitter_AQFP splitterN80ton149n76_( clk_5 , buf_N80_splitterN80ton149n76_1 , 0 , splitterN80ton149n76 );
splitter_AQFP splitterN80ton64n76_( clk_8 , buf_splitterN80ton149n76_splitterN80ton64n76_1 , 0 , splitterN80ton64n76 );
splitter_AQFP splitterN91ton93n345_( clk_3 , buf_N91_splitterN91ton93n345_1 , 0 , splitterN91ton93n345 );
splitter_AQFP splitterN91ton262n345_( clk_5 , splitterN91ton93n345 , 0 , splitterN91ton262n345 );
splitter_AQFP splitterN96ton90n360_( clk_6 , buf_N96_splitterN96ton90n360_1 , 0 , splitterN96ton90n360 );
splitter_AQFP splitterN96ton273n360_( clk_3 , buf_splitterN96ton90n360_splitterN96ton273n360_1 , 0 , splitterN96ton273n360 );
splitter_AQFP splitterfromn61_( clk_5 , n61 , 0 , splitterfromn61 );
splitter_AQFP splitterfromn63_( clk_8 , buf_n63_splitterfromn63_1 , 0 , splitterfromn63 );
splitter_AQFP splittern65ton72N390_( clk_6 , buf_n65_splittern65ton72N390_1 , 0 , splittern65ton72N390 );
splitter_AQFP splittern67ton160n69_( clk_5 , n67 , 0 , splittern67ton160n69 );
splitter_AQFP splitterfromn68_( clk_7 , n68 , 0 , splitterfromn68 );
splitter_AQFP splitterfromn70_( clk_4 , n70 , 0 , splitterfromn70 );
splitter_AQFP splitterfromn71_( clk_6 , buf_n71_splitterfromn71_1 , 0 , splitterfromn71 );
splitter_AQFP splitterfromn73_( clk_6 , n73 , 0 , splitterfromn73 );
splitter_AQFP splitterfromn75_( clk_8 , buf_n75_splitterfromn75_1 , 0 , splitterfromn75 );
splitter_AQFP splitterfromn78_( clk_3 , n78 , 0 , splitterfromn78 );
splitter_AQFP splittern81ton145N447_( clk_6 , n81 , 0 , splittern81ton145N447 );
splitter_AQFP splittern83ton179n88_( clk_7 , n83 , 0 , splittern83ton179n88 );
splitter_AQFP splitterfromn86_( clk_5 , n86 , 0 , splitterfromn86 );
splitter_AQFP splitterfromn92_( clk_3 , n92 , 0 , splitterfromn92 );
splitter_AQFP splitterfromn95_( clk_1 , n95 , 0 , splitterfromn95 );
splitter_AQFP splitterfromn98_( clk_6 , n98 , 0 , splitterfromn98 );
splitter_AQFP splitterfromn101_( clk_3 , n101 , 0 , splitterfromn101 );
splitter_AQFP splitterfromn104_( clk_7 , n104 , 0 , splitterfromn104 );
splitter_AQFP splitterfromn107_( clk_7 , n107 , 0 , splitterfromn107 );
splitter_AQFP splitterfromn110_( clk_3 , n110 , 0 , splitterfromn110 );
splitter_AQFP splitterfromn113_( clk_1 , n113 , 0 , splitterfromn113 );
splitter_AQFP splitterfromn119_( clk_7 , n119 , 0 , splitterfromn119 );
splitter_AQFP splitterfromn122_( clk_5 , n122 , 0 , splitterfromn122 );
splitter_AQFP splitterfromn125_( clk_6 , n125 , 0 , splitterfromn125 );
splitter_AQFP splitterfromn128_( clk_1 , n128 , 0 , splitterfromn128 );
splitter_AQFP splitterfromn131_( clk_6 , n131 , 0 , splitterfromn131 );
splitter_AQFP splitterfromn134_( clk_6 , n134 , 0 , splitterfromn134 );
splitter_AQFP splitterfromn137_( clk_1 , n137 , 0 , splitterfromn137 );
splitter_AQFP splitterfromn140_( clk_6 , n140 , 0 , splitterfromn140 );
splitter_AQFP splitterfromn144_( clk_5 , n144 , 0 , splitterfromn144 );
splitter_AQFP splitterfromn145_( clk_8 , n145 , 0 , splitterfromn145 );
splitter_AQFP splittern147ton148n208_( clk_3 , n147 , 0 , splittern147ton148n208 );
splitter_AQFP splitterfromn150_( clk_8 , n150 , 0 , splitterfromn150 );
splitter_AQFP splittern152ton164n210_( clk_3 , n152 , 0 , splittern152ton164n210 );
splitter_AQFP splittern162ton163n262_( clk_2 , n162 , 0 , splittern162ton163n262 );
splitter_AQFP splittern162ton207n262_( clk_3 , splittern162ton163n262 , 0 , splittern162ton207n262 );
splitter_AQFP splittern162ton273n262_( clk_4 , splittern162ton207n262 , 0 , splittern162ton273n262 );
splitter_AQFP splittern165ton166n175_( clk_6 , n165 , 0 , splittern165ton166n175 );
splitter_AQFP splitterfromn166_( clk_8 , n166 , 0 , splitterfromn166 );
splitter_AQFP splittern167ton168n201_( clk_8 , n167 , 0 , splittern167ton168n201 );
splitter_AQFP splittern168ton169n173_( clk_2 , n168 , 0 , splittern168ton169n173 );
splitter_AQFP splittern179ton253n346_( clk_1 , n179 , 0 , splittern179ton253n346 );
splitter_AQFP splittern179ton315n346_( clk_3 , splittern179ton253n346 , 0 , splittern179ton315n346 );
splitter_AQFP splittern179ton221n346_( clk_5 , splittern179ton315n346 , 0 , splittern179ton221n346 );
splitter_AQFP splittern192ton235n194_( clk_7 , n192 , 0 , splittern192ton235n194 );
splitter_AQFP splittern192ton193n194_( clk_1 , splittern192ton235n194 , 0 , splittern192ton193n194 );
splitter_AQFP splittern193ton228n206_( clk_5 , n193 , 0 , splittern193ton228n206 );
splitter_AQFP splitterfromn194_( clk_5 , n194 , 0 , splitterfromn194 );
splitter_AQFP splittern198ton199n252_( clk_7 , n198 , 0 , splittern198ton199n252 );
splitter_AQFP splittern199ton245n204_( clk_2 , n199 , 0 , splittern199ton245n204 );
splitter_AQFP splitterfromn200_( clk_2 , n200 , 0 , splitterfromn200 );
splitter_AQFP splittern202ton203n247_( clk_3 , n202 , 0 , splittern202ton203n247 );
splitter_AQFP splittern204ton205n230_( clk_6 , n204 , 0 , splittern204ton205n230 );
splitter_AQFP splittern206ton214n297_( clk_1 , n206 , 0 , splittern206ton214n297 );
splitter_AQFP splittern210ton220n212_( clk_8 , n210 , 0 , splittern210ton220n212 );
splitter_AQFP splittern210ton211n212_( clk_2 , splittern210ton220n212 , 0 , splittern210ton211n212 );
splitter_AQFP splittern211ton213n298_( clk_6 , n211 , 0 , splittern211ton213n298 );
splitter_AQFP splitterfromn212_( clk_6 , n212 , 0 , splitterfromn212 );
splitter_AQFP splittern213ton218n215_( clk_8 , n213 , 0 , splittern213ton218n215 );
splitter_AQFP splittern228ton229n233_( clk_7 , n228 , 0 , splittern228ton229n233 );
splitter_AQFP splittern245ton246n250_( clk_4 , n245 , 0 , splittern245ton246n250 );
splitter_AQFP splittern263ton264n282_( clk_2 , n263 , 0 , splittern263ton264n282 );
splitter_AQFP splittern266ton268n292_( clk_2 , n266 , 0 , splittern266ton268n292 );
splitter_AQFP splittern270ton329n272_( clk_1 , n270 , 0 , splittern270ton329n272 );
splitter_AQFP splittern270ton271n272_( clk_3 , splittern270ton329n272 , 0 , splittern270ton271n272 );
splitter_AQFP splittern271ton328n306_( clk_5 , buf_n271_splittern271ton328n306_1 , 0 , splittern271ton328n306 );
splitter_AQFP splitterfromn272_( clk_5 , buf_n272_splitterfromn272_1 , 0 , splitterfromn272 );
splitter_AQFP splittern278ton344n280_( clk_1 , n278 , 0 , splittern278ton344n280 );
splitter_AQFP splittern278ton279n280_( clk_3 , splittern278ton344n280 , 0 , splittern278ton279n280 );
splitter_AQFP splittern279ton343n304_( clk_3 , buf_n279_splittern279ton343n304_1 , 0 , splittern279ton343n304 );
splitter_AQFP splittern279ton337n304_( clk_5 , splittern279ton343n304 , 0 , splittern279ton337n304 );
splitter_AQFP splitterfromn280_( clk_5 , buf_n280_splitterfromn280_1 , 0 , splitterfromn280 );
splitter_AQFP splittern286ton359n288_( clk_1 , n286 , 0 , splittern286ton359n288 );
splitter_AQFP splittern286ton287n288_( clk_3 , splittern286ton359n288 , 0 , splittern286ton287n288 );
splitter_AQFP splittern287ton358n302_( clk_1 , buf_n287_splittern287ton358n302_1 , 0 , splittern287ton358n302 );
splitter_AQFP splittern287ton352n302_( clk_3 , splittern287ton358n302 , 0 , splittern287ton352n302 );
splitter_AQFP splitterfromn288_( clk_2 , buf_n288_splitterfromn288_1 , 0 , splitterfromn288 );
splitter_AQFP splittern294ton314n296_( clk_1 , n294 , 0 , splittern294ton314n296 );
splitter_AQFP splittern294ton295n296_( clk_3 , splittern294ton314n296 , 0 , splittern294ton295n296 );
splitter_AQFP splittern295ton313n300_( clk_8 , buf_n295_splittern295ton313n300_1 , 0 , splittern295ton313n300 );
splitter_AQFP splitterfromn296_( clk_8 , buf_n296_splitterfromn296_1 , 0 , splitterfromn296 );
splitter_AQFP splittern298ton299n312_( clk_4 , n298 , 0 , splittern298ton299n312 );
splitter_AQFP splittern300ton301n354_( clk_7 , n300 , 0 , splittern300ton301n354 );
splitter_AQFP splittern302ton303n339_( clk_2 , n302 , 0 , splittern302ton303n339 );
splitter_AQFP splittern304ton305n324_( clk_5 , n304 , 0 , splittern304ton305n324 );
splitter_AQFP splitterfromn307_( clk_4 , n307 , 0 , splitterfromn307 );
splitter_AQFP splittern322ton327n324_( clk_1 , n322 , 0 , splittern322ton327n324 );
splitter_AQFP splittern322ton323n324_( clk_4 , buf_splittern322ton327n324_splittern322ton323n324_1 , 0 , splittern322ton323n324 );
splitter_AQFP splittern337ton342n339_( clk_1 , n337 , 0 , splittern337ton342n339 );
splitter_AQFP splittern352ton357n354_( clk_6 , n352 , 0 , splittern352ton357n354 );

endmodule