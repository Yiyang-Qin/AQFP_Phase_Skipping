module top( clk_1 , clk_2 , clk_3 , clk_4 , clk_5 , clk_6 , clk_7 , clk_8 , N1 , N101 , N105 , N109 , N113 , N117 , N121 , N125 , N129 , N13 , N130 , N131 , N132 , N133 , N134 , N135 , N136 , N137 , N17 , N21 , N25 , N29 , N33 , N37 , N41 , N45 , N49 , N5 , N53 , N57 , N61 , N65 , N69 , N73 , N77 , N81 , N85 , N89 , N9 , N93 , N97 , N724 , N725 , N726 , N727 , N728 , N729 , N730 , N731 , N732 , N733 , N734 , N735 , N736 , N737 , N738 , N739 , N740 , N741 , N742 , N743 , N744 , N745 , N746 , N747 , N748 , N749 , N750 , N751 , N752 , N753 , N754 , N755 );

input N1 , N101 , N105 , N109 , N113 , N117 , N121 , N125 , N129 , N13 , N130 , N131 , N132 , N133 , N134 , N135 , N136 , N137 , N17 , N21 , N25 , N29 , N33 , N37 , N41 , N45 , N49 , N5 , N53 , N57 , N61 , N65 , N69 , N73 , N77 , N81 , N85 , N89 , N9 , N93 , N97 ;
output N724 , N725 , N726 , N727 , N728 , N729 , N730 , N731 , N732 , N733 , N734 , N735 , N736 , N737 , N738 , N739 , N740 , N741 , N742 , N743 , N744 , N745 , N746 , N747 , N748 , N749 , N750 , N751 , N752 , N753 , N754 , N755 ;
wire n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , buf_N129_n45_1 , buf_N130_n185_1 , buf_N131_n154_1 , buf_N133_n244_1 , buf_N135_n79_2 , buf_N135_n79_1 , buf_n116_splitterfromn116_1 , buf_n154_splitterfromn154_2 , buf_n154_splitterfromn154_1 , buf_n215_splitterfromn215_3 , buf_n215_splitterfromn215_2 , buf_n215_splitterfromn215_1 , buf_splitterN1ton47n284_splitterN1ton283n284_12 , buf_splitterN1ton47n284_splitterN1ton283n284_11 , buf_splitterN1ton47n284_splitterN1ton283n284_10 , buf_splitterN1ton47n284_splitterN1ton283n284_9 , buf_splitterN1ton47n284_splitterN1ton283n284_8 , buf_splitterN1ton47n284_splitterN1ton283n284_7 , buf_splitterN1ton47n284_splitterN1ton283n284_6 , buf_splitterN1ton47n284_splitterN1ton283n284_5 , buf_splitterN1ton47n284_splitterN1ton283n284_4 , buf_splitterN1ton47n284_splitterN1ton283n284_3 , buf_splitterN1ton47n284_splitterN1ton283n284_2 , buf_splitterN1ton47n284_splitterN1ton283n284_1 , buf_splitterN101ton260n402_splitterN101ton401n402_10 , buf_splitterN101ton260n402_splitterN101ton401n402_9 , buf_splitterN101ton260n402_splitterN101ton401n402_8 , buf_splitterN101ton260n402_splitterN101ton401n402_7 , buf_splitterN101ton260n402_splitterN101ton401n402_6 , buf_splitterN101ton260n402_splitterN101ton401n402_5 , buf_splitterN101ton260n402_splitterN101ton401n402_4 , buf_splitterN101ton260n402_splitterN101ton401n402_3 , buf_splitterN101ton260n402_splitterN101ton401n402_2 , buf_splitterN101ton260n402_splitterN101ton401n402_1 , buf_splitterN105ton168n406_splitterN105ton405n406_11 , buf_splitterN105ton168n406_splitterN105ton405n406_10 , buf_splitterN105ton168n406_splitterN105ton405n406_9 , buf_splitterN105ton168n406_splitterN105ton405n406_8 , buf_splitterN105ton168n406_splitterN105ton405n406_7 , buf_splitterN105ton168n406_splitterN105ton405n406_6 , buf_splitterN105ton168n406_splitterN105ton405n406_5 , buf_splitterN105ton168n406_splitterN105ton405n406_4 , buf_splitterN105ton168n406_splitterN105ton405n406_3 , buf_splitterN105ton168n406_splitterN105ton405n406_2 , buf_splitterN105ton168n406_splitterN105ton405n406_1 , buf_splitterN109ton168n410_splitterN109ton409n410_11 , buf_splitterN109ton168n410_splitterN109ton409n410_10 , buf_splitterN109ton168n410_splitterN109ton409n410_9 , buf_splitterN109ton168n410_splitterN109ton409n410_8 , buf_splitterN109ton168n410_splitterN109ton409n410_7 , buf_splitterN109ton168n410_splitterN109ton409n410_6 , buf_splitterN109ton168n410_splitterN109ton409n410_5 , buf_splitterN109ton168n410_splitterN109ton409n410_4 , buf_splitterN109ton168n410_splitterN109ton409n410_3 , buf_splitterN109ton168n410_splitterN109ton409n410_2 , buf_splitterN109ton168n410_splitterN109ton409n410_1 , buf_splitterN113ton241n415_splitterN113ton414n415_10 , buf_splitterN113ton241n415_splitterN113ton414n415_9 , buf_splitterN113ton241n415_splitterN113ton414n415_8 , buf_splitterN113ton241n415_splitterN113ton414n415_7 , buf_splitterN113ton241n415_splitterN113ton414n415_6 , buf_splitterN113ton241n415_splitterN113ton414n415_5 , buf_splitterN113ton241n415_splitterN113ton414n415_4 , buf_splitterN113ton241n415_splitterN113ton414n415_3 , buf_splitterN113ton241n415_splitterN113ton414n415_2 , buf_splitterN113ton241n415_splitterN113ton414n415_1 , buf_splitterN117ton260n419_splitterN117ton418n419_10 , buf_splitterN117ton260n419_splitterN117ton418n419_9 , buf_splitterN117ton260n419_splitterN117ton418n419_8 , buf_splitterN117ton260n419_splitterN117ton418n419_7 , buf_splitterN117ton260n419_splitterN117ton418n419_6 , buf_splitterN117ton260n419_splitterN117ton418n419_5 , buf_splitterN117ton260n419_splitterN117ton418n419_4 , buf_splitterN117ton260n419_splitterN117ton418n419_3 , buf_splitterN117ton260n419_splitterN117ton418n419_2 , buf_splitterN117ton260n419_splitterN117ton418n419_1 , buf_splitterN121ton196n423_splitterN121ton422n423_11 , buf_splitterN121ton196n423_splitterN121ton422n423_10 , buf_splitterN121ton196n423_splitterN121ton422n423_9 , buf_splitterN121ton196n423_splitterN121ton422n423_8 , buf_splitterN121ton196n423_splitterN121ton422n423_7 , buf_splitterN121ton196n423_splitterN121ton422n423_6 , buf_splitterN121ton196n423_splitterN121ton422n423_5 , buf_splitterN121ton196n423_splitterN121ton422n423_4 , buf_splitterN121ton196n423_splitterN121ton422n423_3 , buf_splitterN121ton196n423_splitterN121ton422n423_2 , buf_splitterN121ton196n423_splitterN121ton422n423_1 , buf_splitterN125ton196n427_splitterN125ton426n427_11 , buf_splitterN125ton196n427_splitterN125ton426n427_10 , buf_splitterN125ton196n427_splitterN125ton426n427_9 , buf_splitterN125ton196n427_splitterN125ton426n427_8 , buf_splitterN125ton196n427_splitterN125ton426n427_7 , buf_splitterN125ton196n427_splitterN125ton426n427_6 , buf_splitterN125ton196n427_splitterN125ton426n427_5 , buf_splitterN125ton196n427_splitterN125ton426n427_4 , buf_splitterN125ton196n427_splitterN125ton426n427_3 , buf_splitterN125ton196n427_splitterN125ton426n427_2 , buf_splitterN125ton196n427_splitterN125ton426n427_1 , buf_splitterN13ton219n296_splitterN13ton295n296_11 , buf_splitterN13ton219n296_splitterN13ton295n296_10 , buf_splitterN13ton219n296_splitterN13ton295n296_9 , buf_splitterN13ton219n296_splitterN13ton295n296_8 , buf_splitterN13ton219n296_splitterN13ton295n296_7 , buf_splitterN13ton219n296_splitterN13ton295n296_6 , buf_splitterN13ton219n296_splitterN13ton295n296_5 , buf_splitterN13ton219n296_splitterN13ton295n296_4 , buf_splitterN13ton219n296_splitterN13ton295n296_3 , buf_splitterN13ton219n296_splitterN13ton295n296_2 , buf_splitterN13ton219n296_splitterN13ton295n296_1 , buf_splitterN17ton47n302_splitterN17ton301n302_12 , buf_splitterN17ton47n302_splitterN17ton301n302_11 , buf_splitterN17ton47n302_splitterN17ton301n302_10 , buf_splitterN17ton47n302_splitterN17ton301n302_9 , buf_splitterN17ton47n302_splitterN17ton301n302_8 , buf_splitterN17ton47n302_splitterN17ton301n302_7 , buf_splitterN17ton47n302_splitterN17ton301n302_6 , buf_splitterN17ton47n302_splitterN17ton301n302_5 , buf_splitterN17ton47n302_splitterN17ton301n302_4 , buf_splitterN17ton47n302_splitterN17ton301n302_3 , buf_splitterN17ton47n302_splitterN17ton301n302_2 , buf_splitterN17ton47n302_splitterN17ton301n302_1 , buf_splitterN21ton187n306_splitterN21ton305n306_12 , buf_splitterN21ton187n306_splitterN21ton305n306_11 , buf_splitterN21ton187n306_splitterN21ton305n306_10 , buf_splitterN21ton187n306_splitterN21ton305n306_9 , buf_splitterN21ton187n306_splitterN21ton305n306_8 , buf_splitterN21ton187n306_splitterN21ton305n306_7 , buf_splitterN21ton187n306_splitterN21ton305n306_6 , buf_splitterN21ton187n306_splitterN21ton305n306_5 , buf_splitterN21ton187n306_splitterN21ton305n306_4 , buf_splitterN21ton187n306_splitterN21ton305n306_3 , buf_splitterN21ton187n306_splitterN21ton305n306_2 , buf_splitterN21ton187n306_splitterN21ton305n306_1 , buf_splitterN25ton158n310_splitterN25ton309n310_11 , buf_splitterN25ton158n310_splitterN25ton309n310_10 , buf_splitterN25ton158n310_splitterN25ton309n310_9 , buf_splitterN25ton158n310_splitterN25ton309n310_8 , buf_splitterN25ton158n310_splitterN25ton309n310_7 , buf_splitterN25ton158n310_splitterN25ton309n310_6 , buf_splitterN25ton158n310_splitterN25ton309n310_5 , buf_splitterN25ton158n310_splitterN25ton309n310_4 , buf_splitterN25ton158n310_splitterN25ton309n310_3 , buf_splitterN25ton158n310_splitterN25ton309n310_2 , buf_splitterN25ton158n310_splitterN25ton309n310_1 , buf_splitterN29ton219n314_splitterN29ton313n314_11 , buf_splitterN29ton219n314_splitterN29ton313n314_10 , buf_splitterN29ton219n314_splitterN29ton313n314_9 , buf_splitterN29ton219n314_splitterN29ton313n314_8 , buf_splitterN29ton219n314_splitterN29ton313n314_7 , buf_splitterN29ton219n314_splitterN29ton313n314_6 , buf_splitterN29ton219n314_splitterN29ton313n314_5 , buf_splitterN29ton219n314_splitterN29ton313n314_4 , buf_splitterN29ton219n314_splitterN29ton313n314_3 , buf_splitterN29ton219n314_splitterN29ton313n314_2 , buf_splitterN29ton219n314_splitterN29ton313n314_1 , buf_splitterN33ton42n321_splitterN33ton320n321_11 , buf_splitterN33ton42n321_splitterN33ton320n321_10 , buf_splitterN33ton42n321_splitterN33ton320n321_9 , buf_splitterN33ton42n321_splitterN33ton320n321_8 , buf_splitterN33ton42n321_splitterN33ton320n321_7 , buf_splitterN33ton42n321_splitterN33ton320n321_6 , buf_splitterN33ton42n321_splitterN33ton320n321_5 , buf_splitterN33ton42n321_splitterN33ton320n321_4 , buf_splitterN33ton42n321_splitterN33ton320n321_3 , buf_splitterN33ton42n321_splitterN33ton320n321_2 , buf_splitterN33ton42n321_splitterN33ton320n321_1 , buf_splitterN37ton182n325_splitterN37ton324n325_11 , buf_splitterN37ton182n325_splitterN37ton324n325_10 , buf_splitterN37ton182n325_splitterN37ton324n325_9 , buf_splitterN37ton182n325_splitterN37ton324n325_8 , buf_splitterN37ton182n325_splitterN37ton324n325_7 , buf_splitterN37ton182n325_splitterN37ton324n325_6 , buf_splitterN37ton182n325_splitterN37ton324n325_5 , buf_splitterN37ton182n325_splitterN37ton324n325_4 , buf_splitterN37ton182n325_splitterN37ton324n325_3 , buf_splitterN37ton182n325_splitterN37ton324n325_2 , buf_splitterN37ton182n325_splitterN37ton324n325_1 , buf_splitterN41ton155n329_splitterN41ton328n329_11 , buf_splitterN41ton155n329_splitterN41ton328n329_10 , buf_splitterN41ton155n329_splitterN41ton328n329_9 , buf_splitterN41ton155n329_splitterN41ton328n329_8 , buf_splitterN41ton155n329_splitterN41ton328n329_7 , buf_splitterN41ton155n329_splitterN41ton328n329_6 , buf_splitterN41ton155n329_splitterN41ton328n329_5 , buf_splitterN41ton155n329_splitterN41ton328n329_4 , buf_splitterN41ton155n329_splitterN41ton328n329_3 , buf_splitterN41ton155n329_splitterN41ton328n329_2 , buf_splitterN41ton155n329_splitterN41ton328n329_1 , buf_splitterN45ton216n333_splitterN45ton332n333_11 , buf_splitterN45ton216n333_splitterN45ton332n333_10 , buf_splitterN45ton216n333_splitterN45ton332n333_9 , buf_splitterN45ton216n333_splitterN45ton332n333_8 , buf_splitterN45ton216n333_splitterN45ton332n333_7 , buf_splitterN45ton216n333_splitterN45ton332n333_6 , buf_splitterN45ton216n333_splitterN45ton332n333_5 , buf_splitterN45ton216n333_splitterN45ton332n333_4 , buf_splitterN45ton216n333_splitterN45ton332n333_3 , buf_splitterN45ton216n333_splitterN45ton332n333_2 , buf_splitterN45ton216n333_splitterN45ton332n333_1 , buf_splitterN49ton42n338_splitterN49ton337n338_11 , buf_splitterN49ton42n338_splitterN49ton337n338_10 , buf_splitterN49ton42n338_splitterN49ton337n338_9 , buf_splitterN49ton42n338_splitterN49ton337n338_8 , buf_splitterN49ton42n338_splitterN49ton337n338_7 , buf_splitterN49ton42n338_splitterN49ton337n338_6 , buf_splitterN49ton42n338_splitterN49ton337n338_5 , buf_splitterN49ton42n338_splitterN49ton337n338_4 , buf_splitterN49ton42n338_splitterN49ton337n338_3 , buf_splitterN49ton42n338_splitterN49ton337n338_2 , buf_splitterN49ton42n338_splitterN49ton337n338_1 , buf_splitterN5ton187n288_splitterN5ton287n288_12 , buf_splitterN5ton187n288_splitterN5ton287n288_11 , buf_splitterN5ton187n288_splitterN5ton287n288_10 , buf_splitterN5ton187n288_splitterN5ton287n288_9 , buf_splitterN5ton187n288_splitterN5ton287n288_8 , buf_splitterN5ton187n288_splitterN5ton287n288_7 , buf_splitterN5ton187n288_splitterN5ton287n288_6 , buf_splitterN5ton187n288_splitterN5ton287n288_5 , buf_splitterN5ton187n288_splitterN5ton287n288_4 , buf_splitterN5ton187n288_splitterN5ton287n288_3 , buf_splitterN5ton187n288_splitterN5ton287n288_2 , buf_splitterN5ton187n288_splitterN5ton287n288_1 , buf_splitterN53ton182n342_splitterN53ton341n342_11 , buf_splitterN53ton182n342_splitterN53ton341n342_10 , buf_splitterN53ton182n342_splitterN53ton341n342_9 , buf_splitterN53ton182n342_splitterN53ton341n342_8 , buf_splitterN53ton182n342_splitterN53ton341n342_7 , buf_splitterN53ton182n342_splitterN53ton341n342_6 , buf_splitterN53ton182n342_splitterN53ton341n342_5 , buf_splitterN53ton182n342_splitterN53ton341n342_4 , buf_splitterN53ton182n342_splitterN53ton341n342_3 , buf_splitterN53ton182n342_splitterN53ton341n342_2 , buf_splitterN53ton182n342_splitterN53ton341n342_1 , buf_splitterN57ton155n346_splitterN57ton345n346_11 , buf_splitterN57ton155n346_splitterN57ton345n346_10 , buf_splitterN57ton155n346_splitterN57ton345n346_9 , buf_splitterN57ton155n346_splitterN57ton345n346_8 , buf_splitterN57ton155n346_splitterN57ton345n346_7 , buf_splitterN57ton155n346_splitterN57ton345n346_6 , buf_splitterN57ton155n346_splitterN57ton345n346_5 , buf_splitterN57ton155n346_splitterN57ton345n346_4 , buf_splitterN57ton155n346_splitterN57ton345n346_3 , buf_splitterN57ton155n346_splitterN57ton345n346_2 , buf_splitterN57ton155n346_splitterN57ton345n346_1 , buf_splitterN61ton216n350_splitterN61ton349n350_11 , buf_splitterN61ton216n350_splitterN61ton349n350_10 , buf_splitterN61ton216n350_splitterN61ton349n350_9 , buf_splitterN61ton216n350_splitterN61ton349n350_8 , buf_splitterN61ton216n350_splitterN61ton349n350_7 , buf_splitterN61ton216n350_splitterN61ton349n350_6 , buf_splitterN61ton216n350_splitterN61ton349n350_5 , buf_splitterN61ton216n350_splitterN61ton349n350_4 , buf_splitterN61ton216n350_splitterN61ton349n350_3 , buf_splitterN61ton216n350_splitterN61ton349n350_2 , buf_splitterN61ton216n350_splitterN61ton349n350_1 , buf_splitterN65ton59n363_splitterN65ton362n363_11 , buf_splitterN65ton59n363_splitterN65ton362n363_10 , buf_splitterN65ton59n363_splitterN65ton362n363_9 , buf_splitterN65ton59n363_splitterN65ton362n363_8 , buf_splitterN65ton59n363_splitterN65ton362n363_7 , buf_splitterN65ton59n363_splitterN65ton362n363_6 , buf_splitterN65ton59n363_splitterN65ton362n363_5 , buf_splitterN65ton59n363_splitterN65ton362n363_4 , buf_splitterN65ton59n363_splitterN65ton362n363_3 , buf_splitterN65ton59n363_splitterN65ton362n363_2 , buf_splitterN65ton59n363_splitterN65ton362n363_1 , buf_splitterN69ton59n367_splitterN69ton366n367_11 , buf_splitterN69ton59n367_splitterN69ton366n367_10 , buf_splitterN69ton59n367_splitterN69ton366n367_9 , buf_splitterN69ton59n367_splitterN69ton366n367_8 , buf_splitterN69ton59n367_splitterN69ton366n367_7 , buf_splitterN69ton59n367_splitterN69ton366n367_6 , buf_splitterN69ton59n367_splitterN69ton366n367_5 , buf_splitterN69ton59n367_splitterN69ton366n367_4 , buf_splitterN69ton59n367_splitterN69ton366n367_3 , buf_splitterN69ton59n367_splitterN69ton366n367_2 , buf_splitterN69ton59n367_splitterN69ton366n367_1 , buf_splitterN73ton56n371_splitterN73ton370n371_11 , buf_splitterN73ton56n371_splitterN73ton370n371_10 , buf_splitterN73ton56n371_splitterN73ton370n371_9 , buf_splitterN73ton56n371_splitterN73ton370n371_8 , buf_splitterN73ton56n371_splitterN73ton370n371_7 , buf_splitterN73ton56n371_splitterN73ton370n371_6 , buf_splitterN73ton56n371_splitterN73ton370n371_5 , buf_splitterN73ton56n371_splitterN73ton370n371_4 , buf_splitterN73ton56n371_splitterN73ton370n371_3 , buf_splitterN73ton56n371_splitterN73ton370n371_2 , buf_splitterN73ton56n371_splitterN73ton370n371_1 , buf_splitterN77ton56n375_splitterN77ton374n375_11 , buf_splitterN77ton56n375_splitterN77ton374n375_10 , buf_splitterN77ton56n375_splitterN77ton374n375_9 , buf_splitterN77ton56n375_splitterN77ton374n375_8 , buf_splitterN77ton56n375_splitterN77ton374n375_7 , buf_splitterN77ton56n375_splitterN77ton374n375_6 , buf_splitterN77ton56n375_splitterN77ton374n375_5 , buf_splitterN77ton56n375_splitterN77ton374n375_4 , buf_splitterN77ton56n375_splitterN77ton374n375_3 , buf_splitterN77ton56n375_splitterN77ton374n375_2 , buf_splitterN77ton56n375_splitterN77ton374n375_1 , buf_splitterN81ton68n381_splitterN81ton380n381_11 , buf_splitterN81ton68n381_splitterN81ton380n381_10 , buf_splitterN81ton68n381_splitterN81ton380n381_9 , buf_splitterN81ton68n381_splitterN81ton380n381_8 , buf_splitterN81ton68n381_splitterN81ton380n381_7 , buf_splitterN81ton68n381_splitterN81ton380n381_6 , buf_splitterN81ton68n381_splitterN81ton380n381_5 , buf_splitterN81ton68n381_splitterN81ton380n381_4 , buf_splitterN81ton68n381_splitterN81ton380n381_3 , buf_splitterN81ton68n381_splitterN81ton380n381_2 , buf_splitterN81ton68n381_splitterN81ton380n381_1 , buf_splitterN85ton68n385_splitterN85ton384n385_11 , buf_splitterN85ton68n385_splitterN85ton384n385_10 , buf_splitterN85ton68n385_splitterN85ton384n385_9 , buf_splitterN85ton68n385_splitterN85ton384n385_8 , buf_splitterN85ton68n385_splitterN85ton384n385_7 , buf_splitterN85ton68n385_splitterN85ton384n385_6 , buf_splitterN85ton68n385_splitterN85ton384n385_5 , buf_splitterN85ton68n385_splitterN85ton384n385_4 , buf_splitterN85ton68n385_splitterN85ton384n385_3 , buf_splitterN85ton68n385_splitterN85ton384n385_2 , buf_splitterN85ton68n385_splitterN85ton384n385_1 , buf_splitterN89ton65n389_splitterN89ton388n389_11 , buf_splitterN89ton65n389_splitterN89ton388n389_10 , buf_splitterN89ton65n389_splitterN89ton388n389_9 , buf_splitterN89ton65n389_splitterN89ton388n389_8 , buf_splitterN89ton65n389_splitterN89ton388n389_7 , buf_splitterN89ton65n389_splitterN89ton388n389_6 , buf_splitterN89ton65n389_splitterN89ton388n389_5 , buf_splitterN89ton65n389_splitterN89ton388n389_4 , buf_splitterN89ton65n389_splitterN89ton388n389_3 , buf_splitterN89ton65n389_splitterN89ton388n389_2 , buf_splitterN89ton65n389_splitterN89ton388n389_1 , buf_splitterN9ton158n292_splitterN9ton291n292_11 , buf_splitterN9ton158n292_splitterN9ton291n292_10 , buf_splitterN9ton158n292_splitterN9ton291n292_9 , buf_splitterN9ton158n292_splitterN9ton291n292_8 , buf_splitterN9ton158n292_splitterN9ton291n292_7 , buf_splitterN9ton158n292_splitterN9ton291n292_6 , buf_splitterN9ton158n292_splitterN9ton291n292_5 , buf_splitterN9ton158n292_splitterN9ton291n292_4 , buf_splitterN9ton158n292_splitterN9ton291n292_3 , buf_splitterN9ton158n292_splitterN9ton291n292_2 , buf_splitterN9ton158n292_splitterN9ton291n292_1 , buf_splitterN93ton65n393_splitterN93ton392n393_11 , buf_splitterN93ton65n393_splitterN93ton392n393_10 , buf_splitterN93ton65n393_splitterN93ton392n393_9 , buf_splitterN93ton65n393_splitterN93ton392n393_8 , buf_splitterN93ton65n393_splitterN93ton392n393_7 , buf_splitterN93ton65n393_splitterN93ton392n393_6 , buf_splitterN93ton65n393_splitterN93ton392n393_5 , buf_splitterN93ton65n393_splitterN93ton392n393_4 , buf_splitterN93ton65n393_splitterN93ton392n393_3 , buf_splitterN93ton65n393_splitterN93ton392n393_2 , buf_splitterN93ton65n393_splitterN93ton392n393_1 , buf_splitterN97ton241n398_splitterN97ton397n398_10 , buf_splitterN97ton241n398_splitterN97ton397n398_9 , buf_splitterN97ton241n398_splitterN97ton397n398_8 , buf_splitterN97ton241n398_splitterN97ton397n398_7 , buf_splitterN97ton241n398_splitterN97ton397n398_6 , buf_splitterN97ton241n398_splitterN97ton397n398_5 , buf_splitterN97ton241n398_splitterN97ton397n398_4 , buf_splitterN97ton241n398_splitterN97ton397n398_3 , buf_splitterN97ton241n398_splitterN97ton397n398_2 , buf_splitterN97ton241n398_splitterN97ton397n398_1 , buf_splittern78ton238n336_splittern78ton282n336_4 , buf_splittern78ton238n336_splittern78ton282n336_3 , buf_splittern78ton238n336_splittern78ton282n336_2 , buf_splittern78ton238n336_splittern78ton282n336_1 , buf_splittern115ton353n421_splittern115ton369n421_3 , buf_splittern115ton353n421_splittern115ton369n421_2 , buf_splittern115ton353n421_splittern115ton369n421_1 , buf_splittern152ton353n425_splittern152ton373n425_3 , buf_splittern152ton353n425_splittern152ton373n425_2 , buf_splittern152ton353n425_splittern152ton373n425_1 , buf_splittern153ton355n318_splittern153ton281n318_3 , buf_splittern153ton355n318_splittern153ton281n318_2 , buf_splittern153ton355n318_splittern153ton281n318_1 , buf_splittern181ton236n344_splittern181ton290n344_3 , buf_splittern181ton236n344_splittern181ton290n344_2 , buf_splittern181ton236n344_splittern181ton290n344_1 , buf_splittern209ton210n340_splittern209ton238n340_1 , buf_splittern209ton238n340_splittern209ton286n340_3 , buf_splittern209ton238n340_splittern209ton286n340_2 , buf_splittern209ton238n340_splittern209ton286n340_1 , buf_splitterfromn210_n395_3 , buf_splitterfromn210_n395_2 , buf_splitterfromn210_n395_1 , buf_splitterfromn211_n412_2 , buf_splitterfromn211_n412_1 , buf_splitterfromn212_n360_3 , buf_splitterfromn212_n360_2 , buf_splitterfromn212_n360_1 , buf_splitterfromn213_n378_2 , buf_splitterfromn213_n378_1 , buf_splittern233ton234n348_splittern233ton294n348_2 , buf_splittern233ton234n348_splittern233ton294n348_1 , buf_splitterfromn235_n359_1 , buf_splittern259ton356n413_splittern259ton361n413_3 , buf_splittern259ton356n413_splittern259ton361n413_2 , buf_splittern259ton356n413_splittern259ton361n413_1 , buf_splittern278ton356n417_splittern278ton365n417_3 , buf_splittern278ton356n417_splittern278ton365n417_2 , buf_splittern278ton356n417_splittern278ton365n417_1 , buf_splitterfromn279_n280_3 , buf_splitterfromn279_n280_2 , buf_splitterfromn279_n280_1 , buf_splittern298ton355n335_splittern298ton299n335_3 , buf_splittern298ton355n335_splittern298ton299n335_2 , buf_splittern298ton355n335_splittern298ton299n335_1 , buf_splitterfromn316_n317_3 , buf_splitterfromn316_n317_2 , buf_splitterfromn316_n317_1 , splitterN1ton46n284 , splitterN1ton47n284 , splitterN1ton283n284 , splitterN101ton170n402 , splitterN101ton260n402 , splitterN101ton401n402 , splitterN105ton167n406 , splitterN105ton168n406 , splitterN105ton405n406 , splitterN109ton117n410 , splitterN109ton168n410 , splitterN109ton409n410 , splitterN113ton198n415 , splitterN113ton241n415 , splitterN113ton414n415 , splitterN117ton198n419 , splitterN117ton260n419 , splitterN117ton418n419 , splitterN121ton195n423 , splitterN121ton196n423 , splitterN121ton422n423 , splitterN125ton117n427 , splitterN125ton196n427 , splitterN125ton426n427 , splitterN13ton92n296 , splitterN13ton219n296 , splitterN13ton295n296 , splitterN137ton116n79 , splitterN137ton185n79 , splitterN137ton154n79 , splitterN17ton132n302 , splitterN17ton47n302 , splitterN17ton301n302 , splitterN21ton132n306 , splitterN21ton187n306 , splitterN21ton305n306 , splitterN25ton129n310 , splitterN25ton158n310 , splitterN25ton309n310 , splitterN29ton129n314 , splitterN29ton219n314 , splitterN29ton313n314 , splitterN33ton104n321 , splitterN33ton42n321 , splitterN33ton320n321 , splitterN37ton104n325 , splitterN37ton182n325 , splitterN37ton324n325 , splitterN41ton101n329 , splitterN41ton155n329 , splitterN41ton328n329 , splitterN45ton101n333 , splitterN45ton216n333 , splitterN45ton332n333 , splitterN49ton141n338 , splitterN49ton42n338 , splitterN49ton337n338 , splitterN5ton186n288 , splitterN5ton187n288 , splitterN5ton287n288 , splitterN53ton141n342 , splitterN53ton182n342 , splitterN53ton341n342 , splitterN57ton138n346 , splitterN57ton155n346 , splitterN57ton345n346 , splitterN61ton138n350 , splitterN61ton216n350 , splitterN61ton349n350 , splitterN65ton245n363 , splitterN65ton59n363 , splitterN65ton362n363 , splitterN69ton264n367 , splitterN69ton59n367 , splitterN69ton366n367 , splitterN73ton55n371 , splitterN73ton56n371 , splitterN73ton370n371 , splitterN77ton120n375 , splitterN77ton56n375 , splitterN77ton374n375 , splitterN81ton245n381 , splitterN81ton68n381 , splitterN81ton380n381 , splitterN85ton264n385 , splitterN85ton68n385 , splitterN85ton384n385 , splitterN89ton64n389 , splitterN89ton65n389 , splitterN89ton388n389 , splitterN9ton92n292 , splitterN9ton158n292 , splitterN9ton291n292 , splitterN93ton120n393 , splitterN93ton65n393 , splitterN93ton392n393 , splitterN97ton170n398 , splitterN97ton241n398 , splitterN97ton397n398 , splitterfromn44 , splitterfromn45 , splitterfromn48 , splitterfromn51 , splitterfromn54 , splitterfromn57 , splitterfromn60 , splittern63ton176n74 , splitterfromn66 , splitterfromn69 , splittern72ton73n229 , splitterfromn75 , splittern78ton210n336 , splittern78ton238n336 , splittern78ton282n336 , splitterfromn79 , splitterfromn82 , splitterfromn85 , splitterfromn88 , splitterfromn91 , splitterfromn94 , splitterfromn97 , splittern100ton110n255 , splitterfromn103 , splitterfromn106 , splittern109ton110n274 , splitterfromn112 , splittern115ton153n421 , splittern115ton353n421 , splittern115ton369n421 , splitterfromn116 , splitterfromn119 , splitterfromn122 , splitterfromn125 , splitterfromn128 , splitterfromn131 , splitterfromn134 , splittern137ton147n255 , splitterfromn140 , splitterfromn143 , splittern146ton147n274 , splitterfromn149 , splittern152ton153n425 , splittern152ton353n425 , splittern152ton373n425 , splittern153ton355n318 , splittern153ton281n318 , splitterfromn154 , splitterfromn157 , splitterfromn160 , splitterfromn163 , splitterfromn166 , splitterfromn169 , splitterfromn172 , splittern175ton176n205 , splitterfromn178 , splittern181ton211n344 , splittern181ton236n344 , splittern181ton290n344 , splitterfromn184 , splitterfromn185 , splitterfromn188 , splitterfromn191 , splitterfromn194 , splitterfromn197 , splitterfromn200 , splittern203ton204n229 , splitterfromn206 , splittern209ton210n340 , splittern209ton238n340 , splittern209ton286n340 , splitterfromn210 , splitterfromn211 , splitterfromn212 , splitterfromn213 , splitterfromn215 , splitterfromn218 , splitterfromn221 , splitterfromn224 , splitterfromn227 , splitterfromn230 , splittern233ton235n348 , splittern233ton236n348 , splittern233ton234n348 , splittern233ton294n348 , splitterfromn235 , splitterfromn240 , splitterfromn243 , splitterfromn244 , splitterfromn247 , splitterfromn250 , splitterfromn253 , splitterfromn256 , splittern259ton279n413 , splittern259ton356n413 , splittern259ton361n413 , splitterfromn262 , splitterfromn263 , splitterfromn266 , splitterfromn269 , splitterfromn272 , splitterfromn275 , splittern278ton279n417 , splittern278ton356n417 , splittern278ton365n417 , splitterfromn279 , splitterfromn280 , splittern281ton282n294 , splitterfromn282 , splitterfromn286 , splitterfromn290 , splitterfromn294 , splittern298ton355n335 , splittern298ton299n335 , splittern299ton300n312 , splitterfromn300 , splitterfromn304 , splitterfromn308 , splitterfromn312 , splitterfromn316 , splitterfromn317 , splittern318ton319n331 , splitterfromn319 , splitterfromn323 , splitterfromn327 , splitterfromn331 , splittern335ton336n348 , splitterfromn336 , splitterfromn340 , splitterfromn344 , splitterfromn348 , splitterfromn358 , splitterfromn359 , splittern360ton361n373 , splitterfromn361 , splitterfromn365 , splitterfromn369 , splitterfromn373 , splitterfromn377 , splittern378ton379n391 , splitterfromn379 , splitterfromn383 , splitterfromn387 , splitterfromn391 , splittern395ton396n408 , splitterfromn396 , splitterfromn400 , splitterfromn404 , splitterfromn408 , splittern412ton413n425 , splitterfromn413 , splitterfromn417 , splitterfromn421 , splitterfromn425 ;

PI_AQFP N1_( clk_1 , N1 );
PI_AQFP N101_( clk_1 , N101 );
PI_AQFP N105_( clk_1 , N105 );
PI_AQFP N109_( clk_1 , N109 );
PI_AQFP N113_( clk_1 , N113 );
PI_AQFP N117_( clk_1 , N117 );
PI_AQFP N121_( clk_1 , N121 );
PI_AQFP N125_( clk_1 , N125 );
PI_AQFP N129_( clk_1 , N129 );
PI_AQFP N13_( clk_1 , N13 );
PI_AQFP N130_( clk_1 , N130 );
PI_AQFP N131_( clk_1 , N131 );
PI_AQFP N132_( clk_1 , N132 );
PI_AQFP N133_( clk_1 , N133 );
PI_AQFP N134_( clk_1 , N134 );
PI_AQFP N135_( clk_1 , N135 );
PI_AQFP N136_( clk_1 , N136 );
PI_AQFP N137_( clk_1 , N137 );
PI_AQFP N17_( clk_1 , N17 );
PI_AQFP N21_( clk_1 , N21 );
PI_AQFP N25_( clk_1 , N25 );
PI_AQFP N29_( clk_1 , N29 );
PI_AQFP N33_( clk_1 , N33 );
PI_AQFP N37_( clk_1 , N37 );
PI_AQFP N41_( clk_1 , N41 );
PI_AQFP N45_( clk_1 , N45 );
PI_AQFP N49_( clk_1 , N49 );
PI_AQFP N5_( clk_1 , N5 );
PI_AQFP N53_( clk_1 , N53 );
PI_AQFP N57_( clk_1 , N57 );
PI_AQFP N61_( clk_1 , N61 );
PI_AQFP N65_( clk_1 , N65 );
PI_AQFP N69_( clk_1 , N69 );
PI_AQFP N73_( clk_1 , N73 );
PI_AQFP N77_( clk_1 , N77 );
PI_AQFP N81_( clk_1 , N81 );
PI_AQFP N85_( clk_1 , N85 );
PI_AQFP N89_( clk_1 , N89 );
PI_AQFP N9_( clk_1 , N9 );
PI_AQFP N93_( clk_1 , N93 );
PI_AQFP N97_( clk_1 , N97 );
and_AQFP n42_( clk_6 , splitterN33ton42n321 , splitterN49ton42n338 , 0 , 1 , n42 );
and_AQFP n43_( clk_6 , splitterN33ton42n321 , splitterN49ton42n338 , 1 , 0 , n43 );
or_AQFP n44_( clk_7 , n42 , n43 , 0 , 0 , n44 );
and_AQFP n45_( clk_4 , buf_N129_n45_1 , splitterN137ton185n79 , 0 , 0 , n45 );
and_AQFP n46_( clk_3 , splitterN1ton46n284 , splitterN17ton132n302 , 0 , 1 , n46 );
and_AQFP n47_( clk_4 , splitterN1ton47n284 , splitterN17ton47n302 , 1 , 0 , n47 );
or_AQFP n48_( clk_5 , n46 , n47 , 0 , 0 , n48 );
and_AQFP n49_( clk_7 , splitterfromn45 , splitterfromn48 , 0 , 1 , n49 );
and_AQFP n50_( clk_7 , splitterfromn45 , splitterfromn48 , 1 , 0 , n50 );
or_AQFP n51_( clk_8 , n49 , n50 , 0 , 0 , n51 );
or_AQFP n52_( clk_2 , splitterfromn44 , splitterfromn51 , 0 , 0 , n52 );
and_AQFP n53_( clk_2 , splitterfromn44 , splitterfromn51 , 0 , 0 , n53 );
and_AQFP n54_( clk_3 , n52 , n53 , 0 , 1 , n54 );
or_AQFP n55_( clk_3 , splitterN73ton55n371 , splitterN77ton120n375 , 0 , 0 , n55 );
and_AQFP n56_( clk_4 , splitterN73ton56n371 , splitterN77ton56n375 , 0 , 0 , n56 );
and_AQFP n57_( clk_5 , n55 , n56 , 0 , 1 , n57 );
and_AQFP n58_( clk_3 , splitterN65ton245n363 , splitterN69ton264n367 , 0 , 1 , n58 );
and_AQFP n59_( clk_4 , splitterN65ton59n363 , splitterN69ton59n367 , 1 , 0 , n59 );
or_AQFP n60_( clk_5 , n58 , n59 , 0 , 0 , n60 );
and_AQFP n61_( clk_7 , splitterfromn57 , splitterfromn60 , 1 , 0 , n61 );
and_AQFP n62_( clk_7 , splitterfromn57 , splitterfromn60 , 0 , 1 , n62 );
or_AQFP n63_( clk_8 , n61 , n62 , 0 , 0 , n63 );
or_AQFP n64_( clk_3 , splitterN89ton64n389 , splitterN93ton120n393 , 0 , 0 , n64 );
and_AQFP n65_( clk_4 , splitterN89ton65n389 , splitterN93ton65n393 , 0 , 0 , n65 );
and_AQFP n66_( clk_5 , n64 , n65 , 0 , 1 , n66 );
and_AQFP n67_( clk_3 , splitterN81ton245n381 , splitterN85ton264n385 , 0 , 1 , n67 );
and_AQFP n68_( clk_4 , splitterN81ton68n381 , splitterN85ton68n385 , 1 , 0 , n68 );
or_AQFP n69_( clk_5 , n67 , n68 , 0 , 0 , n69 );
and_AQFP n70_( clk_7 , splitterfromn66 , splitterfromn69 , 1 , 0 , n70 );
and_AQFP n71_( clk_7 , splitterfromn66 , splitterfromn69 , 0 , 1 , n71 );
or_AQFP n72_( clk_8 , n70 , n71 , 0 , 0 , n72 );
and_AQFP n73_( clk_2 , splittern63ton176n74 , splittern72ton73n229 , 0 , 0 , n73 );
or_AQFP n74_( clk_2 , splittern63ton176n74 , splittern72ton73n229 , 0 , 0 , n74 );
and_AQFP n75_( clk_3 , n73 , n74 , 1 , 0 , n75 );
and_AQFP n76_( clk_5 , splitterfromn54 , splitterfromn75 , 1 , 0 , n76 );
and_AQFP n77_( clk_5 , splitterfromn54 , splitterfromn75 , 0 , 1 , n77 );
or_AQFP n78_( clk_6 , n76 , n77 , 0 , 0 , n78 );
and_AQFP n79_( clk_6 , buf_N135_n79_1 , splitterN137ton154n79 , 0 , 0 , n79 );
and_AQFP n80_( clk_3 , splitterN105ton167n406 , splitterN121ton195n423 , 0 , 1 , n80 );
and_AQFP n81_( clk_4 , splitterN105ton168n406 , splitterN121ton196n423 , 1 , 0 , n81 );
or_AQFP n82_( clk_5 , n80 , n81 , 0 , 0 , n82 );
and_AQFP n83_( clk_3 , splitterN73ton55n371 , splitterN89ton64n389 , 0 , 1 , n83 );
and_AQFP n84_( clk_4 , splitterN73ton56n371 , splitterN89ton65n389 , 1 , 0 , n84 );
or_AQFP n85_( clk_5 , n83 , n84 , 0 , 0 , n85 );
and_AQFP n86_( clk_7 , splitterfromn82 , splitterfromn85 , 1 , 0 , n86 );
and_AQFP n87_( clk_7 , splitterfromn82 , splitterfromn85 , 0 , 1 , n87 );
or_AQFP n88_( clk_8 , n86 , n87 , 0 , 0 , n88 );
and_AQFP n89_( clk_2 , splitterfromn79 , splitterfromn88 , 0 , 0 , n89 );
or_AQFP n90_( clk_2 , splitterfromn79 , splitterfromn88 , 0 , 0 , n90 );
and_AQFP n91_( clk_3 , n89 , n90 , 1 , 0 , n91 );
or_AQFP n92_( clk_4 , splitterN13ton92n296 , splitterN9ton92n292 , 0 , 0 , n92 );
and_AQFP n93_( clk_4 , splitterN13ton92n296 , splitterN9ton92n292 , 0 , 0 , n93 );
and_AQFP n94_( clk_5 , n92 , n93 , 0 , 1 , n94 );
and_AQFP n95_( clk_3 , splitterN1ton46n284 , splitterN5ton186n288 , 0 , 1 , n95 );
and_AQFP n96_( clk_4 , splitterN1ton47n284 , splitterN5ton187n288 , 1 , 0 , n96 );
or_AQFP n97_( clk_5 , n95 , n96 , 0 , 0 , n97 );
and_AQFP n98_( clk_7 , splitterfromn94 , splitterfromn97 , 1 , 0 , n98 );
and_AQFP n99_( clk_7 , splitterfromn94 , splitterfromn97 , 0 , 1 , n99 );
or_AQFP n100_( clk_8 , n98 , n99 , 0 , 0 , n100 );
or_AQFP n101_( clk_4 , splitterN41ton101n329 , splitterN45ton101n333 , 0 , 0 , n101 );
and_AQFP n102_( clk_4 , splitterN41ton101n329 , splitterN45ton101n333 , 0 , 0 , n102 );
and_AQFP n103_( clk_5 , n101 , n102 , 0 , 1 , n103 );
and_AQFP n104_( clk_4 , splitterN33ton104n321 , splitterN37ton104n325 , 0 , 1 , n104 );
and_AQFP n105_( clk_4 , splitterN33ton104n321 , splitterN37ton104n325 , 1 , 0 , n105 );
or_AQFP n106_( clk_5 , n104 , n105 , 0 , 0 , n106 );
and_AQFP n107_( clk_7 , splitterfromn103 , splitterfromn106 , 1 , 0 , n107 );
and_AQFP n108_( clk_7 , splitterfromn103 , splitterfromn106 , 0 , 1 , n108 );
or_AQFP n109_( clk_8 , n107 , n108 , 0 , 0 , n109 );
and_AQFP n110_( clk_2 , splittern100ton110n255 , splittern109ton110n274 , 0 , 0 , n110 );
or_AQFP n111_( clk_2 , splittern100ton110n255 , splittern109ton110n274 , 0 , 0 , n111 );
and_AQFP n112_( clk_3 , n110 , n111 , 1 , 0 , n112 );
and_AQFP n113_( clk_5 , splitterfromn91 , splitterfromn112 , 1 , 0 , n113 );
and_AQFP n114_( clk_5 , splitterfromn91 , splitterfromn112 , 0 , 1 , n114 );
or_AQFP n115_( clk_6 , n113 , n114 , 0 , 0 , n115 );
and_AQFP n116_( clk_3 , N136 , splitterN137ton116n79 , 0 , 0 , n116 );
and_AQFP n117_( clk_3 , splitterN109ton117n410 , splitterN125ton117n427 , 0 , 1 , n117 );
and_AQFP n118_( clk_3 , splitterN109ton117n410 , splitterN125ton117n427 , 1 , 0 , n118 );
or_AQFP n119_( clk_4 , n117 , n118 , 0 , 0 , n119 );
and_AQFP n120_( clk_3 , splitterN77ton120n375 , splitterN93ton120n393 , 0 , 1 , n120 );
and_AQFP n121_( clk_3 , splitterN77ton120n375 , splitterN93ton120n393 , 1 , 0 , n121 );
or_AQFP n122_( clk_4 , n120 , n121 , 0 , 0 , n122 );
and_AQFP n123_( clk_6 , splitterfromn119 , splitterfromn122 , 1 , 0 , n123 );
and_AQFP n124_( clk_6 , splitterfromn119 , splitterfromn122 , 0 , 1 , n124 );
or_AQFP n125_( clk_7 , n123 , n124 , 0 , 0 , n125 );
and_AQFP n126_( clk_1 , splitterfromn116 , splitterfromn125 , 0 , 0 , n126 );
or_AQFP n127_( clk_1 , splitterfromn116 , splitterfromn125 , 0 , 0 , n127 );
and_AQFP n128_( clk_2 , n126 , n127 , 1 , 0 , n128 );
or_AQFP n129_( clk_4 , splitterN25ton129n310 , splitterN29ton129n314 , 0 , 0 , n129 );
and_AQFP n130_( clk_4 , splitterN25ton129n310 , splitterN29ton129n314 , 0 , 0 , n130 );
and_AQFP n131_( clk_5 , n129 , n130 , 0 , 1 , n131 );
and_AQFP n132_( clk_3 , splitterN17ton132n302 , splitterN21ton132n306 , 0 , 1 , n132 );
and_AQFP n133_( clk_3 , splitterN17ton132n302 , splitterN21ton132n306 , 1 , 0 , n133 );
or_AQFP n134_( clk_4 , n132 , n133 , 0 , 0 , n134 );
and_AQFP n135_( clk_7 , splitterfromn131 , splitterfromn134 , 1 , 0 , n135 );
and_AQFP n136_( clk_7 , splitterfromn131 , splitterfromn134 , 0 , 1 , n136 );
or_AQFP n137_( clk_8 , n135 , n136 , 0 , 0 , n137 );
or_AQFP n138_( clk_4 , splitterN57ton138n346 , splitterN61ton138n350 , 0 , 0 , n138 );
and_AQFP n139_( clk_4 , splitterN57ton138n346 , splitterN61ton138n350 , 0 , 0 , n139 );
and_AQFP n140_( clk_5 , n138 , n139 , 0 , 1 , n140 );
and_AQFP n141_( clk_4 , splitterN49ton141n338 , splitterN53ton141n342 , 0 , 1 , n141 );
and_AQFP n142_( clk_4 , splitterN49ton141n338 , splitterN53ton141n342 , 1 , 0 , n142 );
or_AQFP n143_( clk_5 , n141 , n142 , 0 , 0 , n143 );
and_AQFP n144_( clk_7 , splitterfromn140 , splitterfromn143 , 1 , 0 , n144 );
and_AQFP n145_( clk_7 , splitterfromn140 , splitterfromn143 , 0 , 1 , n145 );
or_AQFP n146_( clk_8 , n144 , n145 , 0 , 0 , n146 );
and_AQFP n147_( clk_2 , splittern137ton147n255 , splittern146ton147n274 , 0 , 0 , n147 );
or_AQFP n148_( clk_2 , splittern137ton147n255 , splittern146ton147n274 , 0 , 0 , n148 );
and_AQFP n149_( clk_3 , n147 , n148 , 1 , 0 , n149 );
and_AQFP n150_( clk_5 , splitterfromn128 , splitterfromn149 , 1 , 0 , n150 );
and_AQFP n151_( clk_5 , splitterfromn128 , splitterfromn149 , 0 , 1 , n151 );
or_AQFP n152_( clk_6 , n150 , n151 , 0 , 0 , n152 );
and_AQFP n153_( clk_8 , splittern115ton153n421 , splittern152ton153n425 , 0 , 1 , n153 );
and_AQFP n154_( clk_5 , buf_N131_n154_1 , splitterN137ton154n79 , 0 , 0 , n154 );
and_AQFP n155_( clk_6 , splitterN41ton155n329 , splitterN57ton155n346 , 0 , 1 , n155 );
and_AQFP n156_( clk_6 , splitterN41ton155n329 , splitterN57ton155n346 , 1 , 0 , n156 );
or_AQFP n157_( clk_7 , n155 , n156 , 0 , 0 , n157 );
and_AQFP n158_( clk_6 , splitterN25ton158n310 , splitterN9ton158n292 , 1 , 0 , n158 );
and_AQFP n159_( clk_6 , splitterN25ton158n310 , splitterN9ton158n292 , 0 , 1 , n159 );
or_AQFP n160_( clk_7 , n158 , n159 , 0 , 0 , n160 );
and_AQFP n161_( clk_1 , splitterfromn157 , splitterfromn160 , 1 , 0 , n161 );
and_AQFP n162_( clk_1 , splitterfromn157 , splitterfromn160 , 0 , 1 , n162 );
or_AQFP n163_( clk_2 , n161 , n162 , 0 , 0 , n163 );
and_AQFP n164_( clk_4 , splitterfromn154 , splitterfromn163 , 0 , 0 , n164 );
or_AQFP n165_( clk_4 , splitterfromn154 , splitterfromn163 , 0 , 0 , n165 );
and_AQFP n166_( clk_5 , n164 , n165 , 1 , 0 , n166 );
or_AQFP n167_( clk_3 , splitterN105ton167n406 , splitterN109ton117n410 , 0 , 0 , n167 );
and_AQFP n168_( clk_4 , splitterN105ton168n406 , splitterN109ton168n410 , 0 , 0 , n168 );
and_AQFP n169_( clk_5 , n167 , n168 , 0 , 1 , n169 );
and_AQFP n170_( clk_4 , splitterN101ton170n402 , splitterN97ton170n398 , 1 , 0 , n170 );
and_AQFP n171_( clk_4 , splitterN101ton170n402 , splitterN97ton170n398 , 0 , 1 , n171 );
or_AQFP n172_( clk_5 , n170 , n171 , 0 , 0 , n172 );
and_AQFP n173_( clk_7 , splitterfromn169 , splitterfromn172 , 1 , 0 , n173 );
and_AQFP n174_( clk_7 , splitterfromn169 , splitterfromn172 , 0 , 1 , n174 );
or_AQFP n175_( clk_8 , n173 , n174 , 0 , 0 , n175 );
and_AQFP n176_( clk_2 , splittern63ton176n74 , splittern175ton176n205 , 0 , 0 , n176 );
or_AQFP n177_( clk_2 , splittern63ton176n74 , splittern175ton176n205 , 0 , 0 , n177 );
and_AQFP n178_( clk_4 , n176 , n177 , 1 , 0 , n178 );
and_AQFP n179_( clk_7 , splitterfromn166 , splitterfromn178 , 1 , 0 , n179 );
and_AQFP n180_( clk_7 , splitterfromn166 , splitterfromn178 , 0 , 1 , n180 );
or_AQFP n181_( clk_8 , n179 , n180 , 0 , 0 , n181 );
and_AQFP n182_( clk_6 , splitterN37ton182n325 , splitterN53ton182n342 , 0 , 1 , n182 );
and_AQFP n183_( clk_6 , splitterN37ton182n325 , splitterN53ton182n342 , 1 , 0 , n183 );
or_AQFP n184_( clk_8 , n182 , n183 , 0 , 0 , n184 );
and_AQFP n185_( clk_4 , buf_N130_n185_1 , splitterN137ton185n79 , 0 , 0 , n185 );
and_AQFP n186_( clk_3 , splitterN21ton132n306 , splitterN5ton186n288 , 1 , 0 , n186 );
and_AQFP n187_( clk_4 , splitterN21ton187n306 , splitterN5ton187n288 , 0 , 1 , n187 );
or_AQFP n188_( clk_5 , n186 , n187 , 0 , 0 , n188 );
and_AQFP n189_( clk_7 , splitterfromn185 , splitterfromn188 , 0 , 1 , n189 );
and_AQFP n190_( clk_7 , splitterfromn185 , splitterfromn188 , 1 , 0 , n190 );
or_AQFP n191_( clk_8 , n189 , n190 , 0 , 0 , n191 );
or_AQFP n192_( clk_2 , splitterfromn184 , splitterfromn191 , 0 , 0 , n192 );
and_AQFP n193_( clk_2 , splitterfromn184 , splitterfromn191 , 0 , 0 , n193 );
and_AQFP n194_( clk_3 , n192 , n193 , 0 , 1 , n194 );
or_AQFP n195_( clk_3 , splitterN121ton195n423 , splitterN125ton117n427 , 0 , 0 , n195 );
and_AQFP n196_( clk_4 , splitterN121ton196n423 , splitterN125ton196n427 , 0 , 0 , n196 );
and_AQFP n197_( clk_5 , n195 , n196 , 0 , 1 , n197 );
and_AQFP n198_( clk_4 , splitterN113ton198n415 , splitterN117ton198n419 , 0 , 1 , n198 );
and_AQFP n199_( clk_4 , splitterN113ton198n415 , splitterN117ton198n419 , 1 , 0 , n199 );
or_AQFP n200_( clk_5 , n198 , n199 , 0 , 0 , n200 );
and_AQFP n201_( clk_7 , splitterfromn197 , splitterfromn200 , 1 , 0 , n201 );
and_AQFP n202_( clk_7 , splitterfromn197 , splitterfromn200 , 0 , 1 , n202 );
or_AQFP n203_( clk_8 , n201 , n202 , 0 , 0 , n203 );
and_AQFP n204_( clk_2 , splittern175ton176n205 , splittern203ton204n229 , 0 , 0 , n204 );
or_AQFP n205_( clk_2 , splittern175ton176n205 , splittern203ton204n229 , 0 , 0 , n205 );
and_AQFP n206_( clk_3 , n204 , n205 , 1 , 0 , n206 );
and_AQFP n207_( clk_5 , splitterfromn194 , splitterfromn206 , 1 , 0 , n207 );
and_AQFP n208_( clk_5 , splitterfromn194 , splitterfromn206 , 0 , 1 , n208 );
or_AQFP n209_( clk_6 , n207 , n208 , 0 , 0 , n209 );
and_AQFP n210_( clk_8 , splittern78ton210n336 , splittern209ton210n340 , 1 , 0 , n210 );
and_AQFP n211_( clk_2 , splittern181ton211n344 , splitterfromn210 , 1 , 0 , n211 );
and_AQFP n212_( clk_8 , splittern78ton210n336 , splittern209ton210n340 , 0 , 1 , n212 );
and_AQFP n213_( clk_2 , splittern181ton211n344 , splitterfromn212 , 1 , 0 , n213 );
or_AQFP n214_( clk_4 , splitterfromn211 , splitterfromn213 , 0 , 0 , n214 );
and_AQFP n215_( clk_3 , N132 , splitterN137ton116n79 , 0 , 0 , n215 );
and_AQFP n216_( clk_6 , splitterN45ton216n333 , splitterN61ton216n350 , 0 , 1 , n216 );
and_AQFP n217_( clk_6 , splitterN45ton216n333 , splitterN61ton216n350 , 1 , 0 , n217 );
or_AQFP n218_( clk_7 , n216 , n217 , 0 , 0 , n218 );
and_AQFP n219_( clk_6 , splitterN13ton219n296 , splitterN29ton219n314 , 0 , 1 , n219 );
and_AQFP n220_( clk_6 , splitterN13ton219n296 , splitterN29ton219n314 , 1 , 0 , n220 );
or_AQFP n221_( clk_7 , n219 , n220 , 0 , 0 , n221 );
and_AQFP n222_( clk_1 , splitterfromn218 , splitterfromn221 , 1 , 0 , n222 );
and_AQFP n223_( clk_1 , splitterfromn218 , splitterfromn221 , 0 , 1 , n223 );
or_AQFP n224_( clk_2 , n222 , n223 , 0 , 0 , n224 );
and_AQFP n225_( clk_4 , splitterfromn215 , splitterfromn224 , 0 , 0 , n225 );
or_AQFP n226_( clk_4 , splitterfromn215 , splitterfromn224 , 0 , 0 , n226 );
and_AQFP n227_( clk_5 , n225 , n226 , 1 , 0 , n227 );
and_AQFP n228_( clk_3 , splittern72ton73n229 , splittern203ton204n229 , 0 , 0 , n228 );
or_AQFP n229_( clk_3 , splittern72ton73n229 , splittern203ton204n229 , 0 , 0 , n229 );
and_AQFP n230_( clk_4 , n228 , n229 , 1 , 0 , n230 );
and_AQFP n231_( clk_7 , splitterfromn227 , splitterfromn230 , 1 , 0 , n231 );
and_AQFP n232_( clk_7 , splitterfromn227 , splitterfromn230 , 0 , 1 , n232 );
or_AQFP n233_( clk_8 , n231 , n232 , 0 , 0 , n233 );
and_AQFP n234_( clk_5 , n214 , splittern233ton234n348 , 0 , 1 , n234 );
and_AQFP n235_( clk_2 , splittern181ton211n344 , splittern233ton235n348 , 0 , 1 , n235 );
and_AQFP n236_( clk_3 , splittern181ton236n344 , splittern233ton236n348 , 1 , 0 , n236 );
or_AQFP n237_( clk_4 , splitterfromn235 , n236 , 0 , 0 , n237 );
or_AQFP n238_( clk_3 , splittern78ton238n336 , splittern209ton238n340 , 0 , 0 , n238 );
and_AQFP n239_( clk_5 , n237 , n238 , 0 , 1 , n239 );
or_AQFP n240_( clk_6 , n234 , n239 , 0 , 0 , n240 );
and_AQFP n241_( clk_6 , splitterN113ton241n415 , splitterN97ton241n398 , 1 , 0 , n241 );
and_AQFP n242_( clk_6 , splitterN113ton241n415 , splitterN97ton241n398 , 0 , 1 , n242 );
or_AQFP n243_( clk_7 , n241 , n242 , 0 , 0 , n243 );
and_AQFP n244_( clk_4 , buf_N133_n244_1 , splitterN137ton185n79 , 0 , 0 , n244 );
and_AQFP n245_( clk_3 , splitterN65ton245n363 , splitterN81ton245n381 , 0 , 1 , n245 );
and_AQFP n246_( clk_3 , splitterN65ton245n363 , splitterN81ton245n381 , 1 , 0 , n246 );
or_AQFP n247_( clk_4 , n245 , n246 , 0 , 0 , n247 );
and_AQFP n248_( clk_6 , splitterfromn244 , splitterfromn247 , 0 , 1 , n248 );
and_AQFP n249_( clk_6 , splitterfromn244 , splitterfromn247 , 1 , 0 , n249 );
or_AQFP n250_( clk_7 , n248 , n249 , 0 , 0 , n250 );
or_AQFP n251_( clk_1 , splitterfromn243 , splitterfromn250 , 0 , 0 , n251 );
and_AQFP n252_( clk_1 , splitterfromn243 , splitterfromn250 , 0 , 0 , n252 );
and_AQFP n253_( clk_2 , n251 , n252 , 0 , 1 , n253 );
and_AQFP n254_( clk_2 , splittern100ton110n255 , splittern137ton147n255 , 0 , 0 , n254 );
or_AQFP n255_( clk_2 , splittern100ton110n255 , splittern137ton147n255 , 0 , 0 , n255 );
and_AQFP n256_( clk_3 , n254 , n255 , 1 , 0 , n256 );
and_AQFP n257_( clk_5 , splitterfromn253 , splitterfromn256 , 1 , 0 , n257 );
and_AQFP n258_( clk_5 , splitterfromn253 , splitterfromn256 , 0 , 1 , n258 );
or_AQFP n259_( clk_6 , n257 , n258 , 0 , 0 , n259 );
and_AQFP n260_( clk_6 , splitterN101ton260n402 , splitterN117ton260n419 , 0 , 1 , n260 );
and_AQFP n261_( clk_6 , splitterN101ton260n402 , splitterN117ton260n419 , 1 , 0 , n261 );
or_AQFP n262_( clk_7 , n260 , n261 , 0 , 0 , n262 );
and_AQFP n263_( clk_3 , N134 , splitterN137ton116n79 , 0 , 0 , n263 );
and_AQFP n264_( clk_3 , splitterN69ton264n367 , splitterN85ton264n385 , 0 , 1 , n264 );
and_AQFP n265_( clk_3 , splitterN69ton264n367 , splitterN85ton264n385 , 1 , 0 , n265 );
or_AQFP n266_( clk_4 , n264 , n265 , 0 , 0 , n266 );
and_AQFP n267_( clk_6 , splitterfromn263 , splitterfromn266 , 0 , 1 , n267 );
and_AQFP n268_( clk_6 , splitterfromn263 , splitterfromn266 , 1 , 0 , n268 );
or_AQFP n269_( clk_7 , n267 , n268 , 0 , 0 , n269 );
or_AQFP n270_( clk_1 , splitterfromn262 , splitterfromn269 , 0 , 0 , n270 );
and_AQFP n271_( clk_1 , splitterfromn262 , splitterfromn269 , 0 , 0 , n271 );
and_AQFP n272_( clk_2 , n270 , n271 , 0 , 1 , n272 );
and_AQFP n273_( clk_2 , splittern109ton110n274 , splittern146ton147n274 , 0 , 0 , n273 );
or_AQFP n274_( clk_2 , splittern109ton110n274 , splittern146ton147n274 , 0 , 0 , n274 );
and_AQFP n275_( clk_3 , n273 , n274 , 1 , 0 , n275 );
and_AQFP n276_( clk_5 , splitterfromn272 , splitterfromn275 , 1 , 0 , n276 );
and_AQFP n277_( clk_5 , splitterfromn272 , splitterfromn275 , 0 , 1 , n277 );
or_AQFP n278_( clk_6 , n276 , n277 , 0 , 0 , n278 );
and_AQFP n279_( clk_8 , splittern259ton279n413 , splittern278ton279n417 , 0 , 1 , n279 );
and_AQFP n280_( clk_8 , splitterfromn240 , buf_splitterfromn279_n280_1 , 0 , 0 , n280 );
and_AQFP n281_( clk_2 , splittern153ton281n318 , splitterfromn280 , 0 , 0 , n281 );
and_AQFP n282_( clk_4 , splittern78ton282n336 , splittern281ton282n294 , 0 , 0 , n282 );
or_AQFP n283_( clk_6 , splitterN1ton283n284 , splitterfromn282 , 0 , 0 , n283 );
and_AQFP n284_( clk_6 , splitterN1ton283n284 , splitterfromn282 , 0 , 0 , n284 );
and_AQFP n285_( clk_7 , n283 , n284 , 0 , 1 , n285 );
and_AQFP n286_( clk_4 , splittern209ton286n340 , splittern281ton282n294 , 0 , 0 , n286 );
or_AQFP n287_( clk_6 , splitterN5ton287n288 , splitterfromn286 , 0 , 0 , n287 );
and_AQFP n288_( clk_6 , splitterN5ton287n288 , splitterfromn286 , 0 , 0 , n288 );
and_AQFP n289_( clk_7 , n287 , n288 , 0 , 1 , n289 );
and_AQFP n290_( clk_4 , splittern181ton290n344 , splittern281ton282n294 , 0 , 0 , n290 );
and_AQFP n291_( clk_6 , splitterN9ton291n292 , splitterfromn290 , 0 , 0 , n291 );
or_AQFP n292_( clk_6 , splitterN9ton291n292 , splitterfromn290 , 0 , 0 , n292 );
and_AQFP n293_( clk_7 , n291 , n292 , 1 , 0 , n293 );
and_AQFP n294_( clk_4 , splittern233ton294n348 , splittern281ton282n294 , 0 , 0 , n294 );
and_AQFP n295_( clk_6 , splitterN13ton295n296 , splitterfromn294 , 1 , 0 , n295 );
and_AQFP n296_( clk_6 , splitterN13ton295n296 , splitterfromn294 , 0 , 1 , n296 );
or_AQFP n297_( clk_7 , n295 , n296 , 0 , 0 , n297 );
and_AQFP n298_( clk_8 , splittern115ton153n421 , splittern152ton153n425 , 1 , 0 , n298 );
and_AQFP n299_( clk_2 , splitterfromn280 , splittern298ton299n335 , 0 , 0 , n299 );
and_AQFP n300_( clk_4 , splittern78ton282n336 , splittern299ton300n312 , 0 , 0 , n300 );
or_AQFP n301_( clk_6 , splitterN17ton301n302 , splitterfromn300 , 0 , 0 , n301 );
and_AQFP n302_( clk_6 , splitterN17ton301n302 , splitterfromn300 , 0 , 0 , n302 );
and_AQFP n303_( clk_7 , n301 , n302 , 0 , 1 , n303 );
and_AQFP n304_( clk_4 , splittern209ton286n340 , splittern299ton300n312 , 0 , 0 , n304 );
or_AQFP n305_( clk_6 , splitterN21ton305n306 , splitterfromn304 , 0 , 0 , n305 );
and_AQFP n306_( clk_6 , splitterN21ton305n306 , splitterfromn304 , 0 , 0 , n306 );
and_AQFP n307_( clk_7 , n305 , n306 , 0 , 1 , n307 );
and_AQFP n308_( clk_4 , splittern181ton290n344 , splittern299ton300n312 , 0 , 0 , n308 );
and_AQFP n309_( clk_6 , splitterN25ton309n310 , splitterfromn308 , 0 , 0 , n309 );
or_AQFP n310_( clk_6 , splitterN25ton309n310 , splitterfromn308 , 0 , 0 , n310 );
and_AQFP n311_( clk_7 , n309 , n310 , 1 , 0 , n311 );
and_AQFP n312_( clk_4 , splittern233ton294n348 , splittern299ton300n312 , 0 , 0 , n312 );
and_AQFP n313_( clk_6 , splitterN29ton313n314 , splitterfromn312 , 1 , 0 , n313 );
and_AQFP n314_( clk_6 , splitterN29ton313n314 , splitterfromn312 , 0 , 1 , n314 );
or_AQFP n315_( clk_7 , n313 , n314 , 0 , 0 , n315 );
and_AQFP n316_( clk_8 , splittern259ton279n413 , splittern278ton279n417 , 1 , 0 , n316 );
and_AQFP n317_( clk_8 , splitterfromn240 , buf_splitterfromn316_n317_1 , 0 , 0 , n317 );
and_AQFP n318_( clk_2 , splittern153ton281n318 , splitterfromn317 , 0 , 0 , n318 );
and_AQFP n319_( clk_4 , splittern78ton282n336 , splittern318ton319n331 , 0 , 0 , n319 );
or_AQFP n320_( clk_6 , splitterN33ton320n321 , splitterfromn319 , 0 , 0 , n320 );
and_AQFP n321_( clk_6 , splitterN33ton320n321 , splitterfromn319 , 0 , 0 , n321 );
and_AQFP n322_( clk_7 , n320 , n321 , 0 , 1 , n322 );
and_AQFP n323_( clk_4 , splittern209ton286n340 , splittern318ton319n331 , 0 , 0 , n323 );
or_AQFP n324_( clk_6 , splitterN37ton324n325 , splitterfromn323 , 0 , 0 , n324 );
and_AQFP n325_( clk_6 , splitterN37ton324n325 , splitterfromn323 , 0 , 0 , n325 );
and_AQFP n326_( clk_7 , n324 , n325 , 0 , 1 , n326 );
and_AQFP n327_( clk_4 , splittern181ton290n344 , splittern318ton319n331 , 0 , 0 , n327 );
and_AQFP n328_( clk_6 , splitterN41ton328n329 , splitterfromn327 , 0 , 0 , n328 );
or_AQFP n329_( clk_6 , splitterN41ton328n329 , splitterfromn327 , 0 , 0 , n329 );
and_AQFP n330_( clk_7 , n328 , n329 , 1 , 0 , n330 );
and_AQFP n331_( clk_4 , splittern233ton294n348 , splittern318ton319n331 , 0 , 0 , n331 );
or_AQFP n332_( clk_6 , splitterN45ton332n333 , splitterfromn331 , 0 , 0 , n332 );
and_AQFP n333_( clk_6 , splitterN45ton332n333 , splitterfromn331 , 0 , 0 , n333 );
and_AQFP n334_( clk_7 , n332 , n333 , 0 , 1 , n334 );
and_AQFP n335_( clk_2 , splittern298ton299n335 , splitterfromn317 , 0 , 0 , n335 );
and_AQFP n336_( clk_4 , splittern78ton282n336 , splittern335ton336n348 , 0 , 0 , n336 );
or_AQFP n337_( clk_6 , splitterN49ton337n338 , splitterfromn336 , 0 , 0 , n337 );
and_AQFP n338_( clk_6 , splitterN49ton337n338 , splitterfromn336 , 0 , 0 , n338 );
and_AQFP n339_( clk_7 , n337 , n338 , 0 , 1 , n339 );
and_AQFP n340_( clk_4 , splittern209ton286n340 , splittern335ton336n348 , 0 , 0 , n340 );
or_AQFP n341_( clk_6 , splitterN53ton341n342 , splitterfromn340 , 0 , 0 , n341 );
and_AQFP n342_( clk_6 , splitterN53ton341n342 , splitterfromn340 , 0 , 0 , n342 );
and_AQFP n343_( clk_7 , n341 , n342 , 0 , 1 , n343 );
and_AQFP n344_( clk_4 , splittern181ton290n344 , splittern335ton336n348 , 0 , 0 , n344 );
and_AQFP n345_( clk_6 , splitterN57ton345n346 , splitterfromn344 , 0 , 0 , n345 );
or_AQFP n346_( clk_6 , splitterN57ton345n346 , splitterfromn344 , 0 , 0 , n346 );
and_AQFP n347_( clk_7 , n345 , n346 , 1 , 0 , n347 );
and_AQFP n348_( clk_4 , splittern233ton294n348 , splittern335ton336n348 , 0 , 0 , n348 );
and_AQFP n349_( clk_6 , splitterN61ton349n350 , splitterfromn348 , 0 , 0 , n349 );
or_AQFP n350_( clk_6 , splitterN61ton349n350 , splitterfromn348 , 0 , 0 , n350 );
and_AQFP n351_( clk_7 , n349 , n350 , 1 , 0 , n351 );
or_AQFP n352_( clk_2 , splitterfromn279 , splitterfromn316 , 0 , 0 , n352 );
or_AQFP n353_( clk_2 , splittern115ton353n421 , splittern152ton353n425 , 0 , 0 , n353 );
and_AQFP n354_( clk_3 , n352 , n353 , 0 , 1 , n354 );
or_AQFP n355_( clk_2 , splittern153ton355n318 , splittern298ton355n335 , 0 , 0 , n355 );
or_AQFP n356_( clk_2 , splittern259ton356n413 , splittern278ton356n417 , 0 , 0 , n356 );
and_AQFP n357_( clk_3 , n355 , n356 , 0 , 1 , n357 );
or_AQFP n358_( clk_4 , n354 , n357 , 0 , 0 , n358 );
and_AQFP n359_( clk_6 , buf_splitterfromn235_n359_1 , splitterfromn358 , 0 , 0 , n359 );
and_AQFP n360_( clk_8 , buf_splitterfromn212_n360_1 , splitterfromn359 , 0 , 0 , n360 );
and_AQFP n361_( clk_2 , splittern259ton361n413 , splittern360ton361n373 , 0 , 0 , n361 );
or_AQFP n362_( clk_4 , splitterN65ton362n363 , splitterfromn361 , 0 , 0 , n362 );
and_AQFP n363_( clk_4 , splitterN65ton362n363 , splitterfromn361 , 0 , 0 , n363 );
and_AQFP n364_( clk_6 , n362 , n363 , 0 , 1 , n364 );
and_AQFP n365_( clk_2 , splittern278ton365n417 , splittern360ton361n373 , 0 , 0 , n365 );
or_AQFP n366_( clk_4 , splitterN69ton366n367 , splitterfromn365 , 0 , 0 , n366 );
and_AQFP n367_( clk_4 , splitterN69ton366n367 , splitterfromn365 , 0 , 0 , n367 );
and_AQFP n368_( clk_6 , n366 , n367 , 0 , 1 , n368 );
and_AQFP n369_( clk_2 , splittern115ton369n421 , splittern360ton361n373 , 0 , 0 , n369 );
and_AQFP n370_( clk_4 , splitterN73ton370n371 , splitterfromn369 , 1 , 0 , n370 );
and_AQFP n371_( clk_4 , splitterN73ton370n371 , splitterfromn369 , 0 , 1 , n371 );
or_AQFP n372_( clk_6 , n370 , n371 , 0 , 0 , n372 );
and_AQFP n373_( clk_2 , splittern152ton373n425 , splittern360ton361n373 , 0 , 0 , n373 );
and_AQFP n374_( clk_4 , splitterN77ton374n375 , splitterfromn373 , 0 , 0 , n374 );
or_AQFP n375_( clk_4 , splitterN77ton374n375 , splitterfromn373 , 0 , 0 , n375 );
and_AQFP n376_( clk_6 , n374 , n375 , 1 , 0 , n376 );
and_AQFP n377_( clk_6 , splittern233ton234n348 , splitterfromn358 , 0 , 0 , n377 );
and_AQFP n378_( clk_8 , buf_splitterfromn213_n378_1 , splitterfromn377 , 0 , 0 , n378 );
and_AQFP n379_( clk_2 , splittern259ton361n413 , splittern378ton379n391 , 0 , 0 , n379 );
or_AQFP n380_( clk_4 , splitterN81ton380n381 , splitterfromn379 , 0 , 0 , n380 );
and_AQFP n381_( clk_4 , splitterN81ton380n381 , splitterfromn379 , 0 , 0 , n381 );
and_AQFP n382_( clk_6 , n380 , n381 , 0 , 1 , n382 );
and_AQFP n383_( clk_2 , splittern278ton365n417 , splittern378ton379n391 , 0 , 0 , n383 );
or_AQFP n384_( clk_4 , splitterN85ton384n385 , splitterfromn383 , 0 , 0 , n384 );
and_AQFP n385_( clk_4 , splitterN85ton384n385 , splitterfromn383 , 0 , 0 , n385 );
and_AQFP n386_( clk_6 , n384 , n385 , 0 , 1 , n386 );
and_AQFP n387_( clk_2 , splittern115ton369n421 , splittern378ton379n391 , 0 , 0 , n387 );
and_AQFP n388_( clk_4 , splitterN89ton388n389 , splitterfromn387 , 0 , 0 , n388 );
or_AQFP n389_( clk_4 , splitterN89ton388n389 , splitterfromn387 , 0 , 0 , n389 );
and_AQFP n390_( clk_6 , n388 , n389 , 1 , 0 , n390 );
and_AQFP n391_( clk_2 , splittern152ton373n425 , splittern378ton379n391 , 0 , 0 , n391 );
or_AQFP n392_( clk_4 , splitterN93ton392n393 , splitterfromn391 , 0 , 0 , n392 );
and_AQFP n393_( clk_4 , splitterN93ton392n393 , splitterfromn391 , 0 , 0 , n393 );
and_AQFP n394_( clk_6 , n392 , n393 , 0 , 1 , n394 );
and_AQFP n395_( clk_8 , buf_splitterfromn210_n395_1 , splitterfromn359 , 0 , 0 , n395 );
and_AQFP n396_( clk_2 , splittern259ton361n413 , splittern395ton396n408 , 0 , 0 , n396 );
or_AQFP n397_( clk_4 , splitterN97ton397n398 , splitterfromn396 , 0 , 0 , n397 );
and_AQFP n398_( clk_4 , splitterN97ton397n398 , splitterfromn396 , 0 , 0 , n398 );
and_AQFP n399_( clk_6 , n397 , n398 , 0 , 1 , n399 );
and_AQFP n400_( clk_2 , splittern278ton365n417 , splittern395ton396n408 , 0 , 0 , n400 );
or_AQFP n401_( clk_4 , splitterN101ton401n402 , splitterfromn400 , 0 , 0 , n401 );
and_AQFP n402_( clk_4 , splitterN101ton401n402 , splitterfromn400 , 0 , 0 , n402 );
and_AQFP n403_( clk_6 , n401 , n402 , 0 , 1 , n403 );
and_AQFP n404_( clk_2 , splittern115ton369n421 , splittern395ton396n408 , 0 , 0 , n404 );
and_AQFP n405_( clk_4 , splitterN105ton405n406 , splitterfromn404 , 1 , 0 , n405 );
and_AQFP n406_( clk_4 , splitterN105ton405n406 , splitterfromn404 , 0 , 1 , n406 );
or_AQFP n407_( clk_6 , n405 , n406 , 0 , 0 , n407 );
and_AQFP n408_( clk_2 , splittern152ton373n425 , splittern395ton396n408 , 0 , 0 , n408 );
and_AQFP n409_( clk_4 , splitterN109ton409n410 , splitterfromn408 , 0 , 0 , n409 );
or_AQFP n410_( clk_4 , splitterN109ton409n410 , splitterfromn408 , 0 , 0 , n410 );
and_AQFP n411_( clk_6 , n409 , n410 , 1 , 0 , n411 );
and_AQFP n412_( clk_8 , buf_splitterfromn211_n412_1 , splitterfromn377 , 0 , 0 , n412 );
and_AQFP n413_( clk_2 , splittern259ton361n413 , splittern412ton413n425 , 0 , 0 , n413 );
or_AQFP n414_( clk_4 , splitterN113ton414n415 , splitterfromn413 , 0 , 0 , n414 );
and_AQFP n415_( clk_4 , splitterN113ton414n415 , splitterfromn413 , 0 , 0 , n415 );
and_AQFP n416_( clk_6 , n414 , n415 , 0 , 1 , n416 );
and_AQFP n417_( clk_2 , splittern278ton365n417 , splittern412ton413n425 , 0 , 0 , n417 );
or_AQFP n418_( clk_4 , splitterN117ton418n419 , splitterfromn417 , 0 , 0 , n418 );
and_AQFP n419_( clk_4 , splitterN117ton418n419 , splitterfromn417 , 0 , 0 , n419 );
and_AQFP n420_( clk_6 , n418 , n419 , 0 , 1 , n420 );
and_AQFP n421_( clk_2 , splittern115ton369n421 , splittern412ton413n425 , 0 , 0 , n421 );
and_AQFP n422_( clk_4 , splitterN121ton422n423 , splitterfromn421 , 0 , 0 , n422 );
or_AQFP n423_( clk_4 , splitterN121ton422n423 , splitterfromn421 , 0 , 0 , n423 );
and_AQFP n424_( clk_6 , n422 , n423 , 1 , 0 , n424 );
and_AQFP n425_( clk_2 , splittern152ton373n425 , splittern412ton413n425 , 0 , 0 , n425 );
or_AQFP n426_( clk_4 , splitterN125ton426n427 , splitterfromn425 , 0 , 0 , n426 );
and_AQFP n427_( clk_4 , splitterN125ton426n427 , splitterfromn425 , 0 , 0 , n427 );
and_AQFP n428_( clk_6 , n426 , n427 , 0 , 1 , n428 );
PO_AQFP N724_( clk_8 , n285 , 0 , N724 );
PO_AQFP N725_( clk_8 , n289 , 0 , N725 );
PO_AQFP N726_( clk_8 , n293 , 0 , N726 );
PO_AQFP N727_( clk_8 , n297 , 0 , N727 );
PO_AQFP N728_( clk_8 , n303 , 0 , N728 );
PO_AQFP N729_( clk_8 , n307 , 0 , N729 );
PO_AQFP N730_( clk_8 , n311 , 0 , N730 );
PO_AQFP N731_( clk_8 , n315 , 0 , N731 );
PO_AQFP N732_( clk_8 , n322 , 0 , N732 );
PO_AQFP N733_( clk_8 , n326 , 0 , N733 );
PO_AQFP N734_( clk_8 , n330 , 0 , N734 );
PO_AQFP N735_( clk_8 , n334 , 0 , N735 );
PO_AQFP N736_( clk_8 , n339 , 0 , N736 );
PO_AQFP N737_( clk_8 , n343 , 0 , N737 );
PO_AQFP N738_( clk_8 , n347 , 0 , N738 );
PO_AQFP N739_( clk_8 , n351 , 0 , N739 );
PO_AQFP N740_( clk_8 , n364 , 0 , N740 );
PO_AQFP N741_( clk_8 , n368 , 0 , N741 );
PO_AQFP N742_( clk_8 , n372 , 0 , N742 );
PO_AQFP N743_( clk_8 , n376 , 0 , N743 );
PO_AQFP N744_( clk_8 , n382 , 0 , N744 );
PO_AQFP N745_( clk_8 , n386 , 0 , N745 );
PO_AQFP N746_( clk_8 , n390 , 0 , N746 );
PO_AQFP N747_( clk_8 , n394 , 0 , N747 );
PO_AQFP N748_( clk_8 , n399 , 0 , N748 );
PO_AQFP N749_( clk_8 , n403 , 0 , N749 );
PO_AQFP N750_( clk_8 , n407 , 0 , N750 );
PO_AQFP N751_( clk_8 , n411 , 0 , N751 );
PO_AQFP N752_( clk_8 , n416 , 0 , N752 );
PO_AQFP N753_( clk_8 , n420 , 0 , N753 );
PO_AQFP N754_( clk_8 , n424 , 0 , N754 );
PO_AQFP N755_( clk_8 , n428 , 0 , N755 );
buf_AQFP buf_N129_n45_1_( clk_3 , N129 , 0 , buf_N129_n45_1 );
buf_AQFP buf_N130_n185_1_( clk_3 , N130 , 0 , buf_N130_n185_1 );
buf_AQFP buf_N131_n154_1_( clk_3 , N131 , 0 , buf_N131_n154_1 );
buf_AQFP buf_N133_n244_1_( clk_3 , N133 , 0 , buf_N133_n244_1 );
buf_AQFP buf_N135_n79_2_( clk_3 , N135 , 0 , buf_N135_n79_2 );
buf_AQFP buf_N135_n79_1_( clk_5 , buf_N135_n79_2 , 0 , buf_N135_n79_1 );
buf_AQFP buf_n116_splitterfromn116_1_( clk_5 , n116 , 0 , buf_n116_splitterfromn116_1 );
buf_AQFP buf_n154_splitterfromn154_2_( clk_7 , n154 , 0 , buf_n154_splitterfromn154_2 );
buf_AQFP buf_n154_splitterfromn154_1_( clk_1 , buf_n154_splitterfromn154_2 , 0 , buf_n154_splitterfromn154_1 );
buf_AQFP buf_n215_splitterfromn215_3_( clk_5 , n215 , 0 , buf_n215_splitterfromn215_3 );
buf_AQFP buf_n215_splitterfromn215_2_( clk_7 , buf_n215_splitterfromn215_3 , 0 , buf_n215_splitterfromn215_2 );
buf_AQFP buf_n215_splitterfromn215_1_( clk_1 , buf_n215_splitterfromn215_2 , 0 , buf_n215_splitterfromn215_1 );
buf_AQFP buf_splitterN1ton47n284_splitterN1ton283n284_12_( clk_5 , splitterN1ton47n284 , 0 , buf_splitterN1ton47n284_splitterN1ton283n284_12 );
buf_AQFP buf_splitterN1ton47n284_splitterN1ton283n284_11_( clk_7 , buf_splitterN1ton47n284_splitterN1ton283n284_12 , 0 , buf_splitterN1ton47n284_splitterN1ton283n284_11 );
buf_AQFP buf_splitterN1ton47n284_splitterN1ton283n284_10_( clk_1 , buf_splitterN1ton47n284_splitterN1ton283n284_11 , 0 , buf_splitterN1ton47n284_splitterN1ton283n284_10 );
buf_AQFP buf_splitterN1ton47n284_splitterN1ton283n284_9_( clk_3 , buf_splitterN1ton47n284_splitterN1ton283n284_10 , 0 , buf_splitterN1ton47n284_splitterN1ton283n284_9 );
buf_AQFP buf_splitterN1ton47n284_splitterN1ton283n284_8_( clk_5 , buf_splitterN1ton47n284_splitterN1ton283n284_9 , 0 , buf_splitterN1ton47n284_splitterN1ton283n284_8 );
buf_AQFP buf_splitterN1ton47n284_splitterN1ton283n284_7_( clk_7 , buf_splitterN1ton47n284_splitterN1ton283n284_8 , 0 , buf_splitterN1ton47n284_splitterN1ton283n284_7 );
buf_AQFP buf_splitterN1ton47n284_splitterN1ton283n284_6_( clk_1 , buf_splitterN1ton47n284_splitterN1ton283n284_7 , 0 , buf_splitterN1ton47n284_splitterN1ton283n284_6 );
buf_AQFP buf_splitterN1ton47n284_splitterN1ton283n284_5_( clk_3 , buf_splitterN1ton47n284_splitterN1ton283n284_6 , 0 , buf_splitterN1ton47n284_splitterN1ton283n284_5 );
buf_AQFP buf_splitterN1ton47n284_splitterN1ton283n284_4_( clk_5 , buf_splitterN1ton47n284_splitterN1ton283n284_5 , 0 , buf_splitterN1ton47n284_splitterN1ton283n284_4 );
buf_AQFP buf_splitterN1ton47n284_splitterN1ton283n284_3_( clk_7 , buf_splitterN1ton47n284_splitterN1ton283n284_4 , 0 , buf_splitterN1ton47n284_splitterN1ton283n284_3 );
buf_AQFP buf_splitterN1ton47n284_splitterN1ton283n284_2_( clk_1 , buf_splitterN1ton47n284_splitterN1ton283n284_3 , 0 , buf_splitterN1ton47n284_splitterN1ton283n284_2 );
buf_AQFP buf_splitterN1ton47n284_splitterN1ton283n284_1_( clk_3 , buf_splitterN1ton47n284_splitterN1ton283n284_2 , 0 , buf_splitterN1ton47n284_splitterN1ton283n284_1 );
buf_AQFP buf_splitterN101ton260n402_splitterN101ton401n402_10_( clk_7 , splitterN101ton260n402 , 0 , buf_splitterN101ton260n402_splitterN101ton401n402_10 );
buf_AQFP buf_splitterN101ton260n402_splitterN101ton401n402_9_( clk_1 , buf_splitterN101ton260n402_splitterN101ton401n402_10 , 0 , buf_splitterN101ton260n402_splitterN101ton401n402_9 );
buf_AQFP buf_splitterN101ton260n402_splitterN101ton401n402_8_( clk_3 , buf_splitterN101ton260n402_splitterN101ton401n402_9 , 0 , buf_splitterN101ton260n402_splitterN101ton401n402_8 );
buf_AQFP buf_splitterN101ton260n402_splitterN101ton401n402_7_( clk_5 , buf_splitterN101ton260n402_splitterN101ton401n402_8 , 0 , buf_splitterN101ton260n402_splitterN101ton401n402_7 );
buf_AQFP buf_splitterN101ton260n402_splitterN101ton401n402_6_( clk_7 , buf_splitterN101ton260n402_splitterN101ton401n402_7 , 0 , buf_splitterN101ton260n402_splitterN101ton401n402_6 );
buf_AQFP buf_splitterN101ton260n402_splitterN101ton401n402_5_( clk_1 , buf_splitterN101ton260n402_splitterN101ton401n402_6 , 0 , buf_splitterN101ton260n402_splitterN101ton401n402_5 );
buf_AQFP buf_splitterN101ton260n402_splitterN101ton401n402_4_( clk_3 , buf_splitterN101ton260n402_splitterN101ton401n402_5 , 0 , buf_splitterN101ton260n402_splitterN101ton401n402_4 );
buf_AQFP buf_splitterN101ton260n402_splitterN101ton401n402_3_( clk_5 , buf_splitterN101ton260n402_splitterN101ton401n402_4 , 0 , buf_splitterN101ton260n402_splitterN101ton401n402_3 );
buf_AQFP buf_splitterN101ton260n402_splitterN101ton401n402_2_( clk_7 , buf_splitterN101ton260n402_splitterN101ton401n402_3 , 0 , buf_splitterN101ton260n402_splitterN101ton401n402_2 );
buf_AQFP buf_splitterN101ton260n402_splitterN101ton401n402_1_( clk_1 , buf_splitterN101ton260n402_splitterN101ton401n402_2 , 0 , buf_splitterN101ton260n402_splitterN101ton401n402_1 );
buf_AQFP buf_splitterN105ton168n406_splitterN105ton405n406_11_( clk_5 , splitterN105ton168n406 , 0 , buf_splitterN105ton168n406_splitterN105ton405n406_11 );
buf_AQFP buf_splitterN105ton168n406_splitterN105ton405n406_10_( clk_7 , buf_splitterN105ton168n406_splitterN105ton405n406_11 , 0 , buf_splitterN105ton168n406_splitterN105ton405n406_10 );
buf_AQFP buf_splitterN105ton168n406_splitterN105ton405n406_9_( clk_1 , buf_splitterN105ton168n406_splitterN105ton405n406_10 , 0 , buf_splitterN105ton168n406_splitterN105ton405n406_9 );
buf_AQFP buf_splitterN105ton168n406_splitterN105ton405n406_8_( clk_3 , buf_splitterN105ton168n406_splitterN105ton405n406_9 , 0 , buf_splitterN105ton168n406_splitterN105ton405n406_8 );
buf_AQFP buf_splitterN105ton168n406_splitterN105ton405n406_7_( clk_5 , buf_splitterN105ton168n406_splitterN105ton405n406_8 , 0 , buf_splitterN105ton168n406_splitterN105ton405n406_7 );
buf_AQFP buf_splitterN105ton168n406_splitterN105ton405n406_6_( clk_7 , buf_splitterN105ton168n406_splitterN105ton405n406_7 , 0 , buf_splitterN105ton168n406_splitterN105ton405n406_6 );
buf_AQFP buf_splitterN105ton168n406_splitterN105ton405n406_5_( clk_1 , buf_splitterN105ton168n406_splitterN105ton405n406_6 , 0 , buf_splitterN105ton168n406_splitterN105ton405n406_5 );
buf_AQFP buf_splitterN105ton168n406_splitterN105ton405n406_4_( clk_3 , buf_splitterN105ton168n406_splitterN105ton405n406_5 , 0 , buf_splitterN105ton168n406_splitterN105ton405n406_4 );
buf_AQFP buf_splitterN105ton168n406_splitterN105ton405n406_3_( clk_5 , buf_splitterN105ton168n406_splitterN105ton405n406_4 , 0 , buf_splitterN105ton168n406_splitterN105ton405n406_3 );
buf_AQFP buf_splitterN105ton168n406_splitterN105ton405n406_2_( clk_7 , buf_splitterN105ton168n406_splitterN105ton405n406_3 , 0 , buf_splitterN105ton168n406_splitterN105ton405n406_2 );
buf_AQFP buf_splitterN105ton168n406_splitterN105ton405n406_1_( clk_1 , buf_splitterN105ton168n406_splitterN105ton405n406_2 , 0 , buf_splitterN105ton168n406_splitterN105ton405n406_1 );
buf_AQFP buf_splitterN109ton168n410_splitterN109ton409n410_11_( clk_5 , splitterN109ton168n410 , 0 , buf_splitterN109ton168n410_splitterN109ton409n410_11 );
buf_AQFP buf_splitterN109ton168n410_splitterN109ton409n410_10_( clk_7 , buf_splitterN109ton168n410_splitterN109ton409n410_11 , 0 , buf_splitterN109ton168n410_splitterN109ton409n410_10 );
buf_AQFP buf_splitterN109ton168n410_splitterN109ton409n410_9_( clk_1 , buf_splitterN109ton168n410_splitterN109ton409n410_10 , 0 , buf_splitterN109ton168n410_splitterN109ton409n410_9 );
buf_AQFP buf_splitterN109ton168n410_splitterN109ton409n410_8_( clk_3 , buf_splitterN109ton168n410_splitterN109ton409n410_9 , 0 , buf_splitterN109ton168n410_splitterN109ton409n410_8 );
buf_AQFP buf_splitterN109ton168n410_splitterN109ton409n410_7_( clk_5 , buf_splitterN109ton168n410_splitterN109ton409n410_8 , 0 , buf_splitterN109ton168n410_splitterN109ton409n410_7 );
buf_AQFP buf_splitterN109ton168n410_splitterN109ton409n410_6_( clk_7 , buf_splitterN109ton168n410_splitterN109ton409n410_7 , 0 , buf_splitterN109ton168n410_splitterN109ton409n410_6 );
buf_AQFP buf_splitterN109ton168n410_splitterN109ton409n410_5_( clk_1 , buf_splitterN109ton168n410_splitterN109ton409n410_6 , 0 , buf_splitterN109ton168n410_splitterN109ton409n410_5 );
buf_AQFP buf_splitterN109ton168n410_splitterN109ton409n410_4_( clk_3 , buf_splitterN109ton168n410_splitterN109ton409n410_5 , 0 , buf_splitterN109ton168n410_splitterN109ton409n410_4 );
buf_AQFP buf_splitterN109ton168n410_splitterN109ton409n410_3_( clk_5 , buf_splitterN109ton168n410_splitterN109ton409n410_4 , 0 , buf_splitterN109ton168n410_splitterN109ton409n410_3 );
buf_AQFP buf_splitterN109ton168n410_splitterN109ton409n410_2_( clk_7 , buf_splitterN109ton168n410_splitterN109ton409n410_3 , 0 , buf_splitterN109ton168n410_splitterN109ton409n410_2 );
buf_AQFP buf_splitterN109ton168n410_splitterN109ton409n410_1_( clk_1 , buf_splitterN109ton168n410_splitterN109ton409n410_2 , 0 , buf_splitterN109ton168n410_splitterN109ton409n410_1 );
buf_AQFP buf_splitterN113ton241n415_splitterN113ton414n415_10_( clk_7 , splitterN113ton241n415 , 0 , buf_splitterN113ton241n415_splitterN113ton414n415_10 );
buf_AQFP buf_splitterN113ton241n415_splitterN113ton414n415_9_( clk_1 , buf_splitterN113ton241n415_splitterN113ton414n415_10 , 0 , buf_splitterN113ton241n415_splitterN113ton414n415_9 );
buf_AQFP buf_splitterN113ton241n415_splitterN113ton414n415_8_( clk_3 , buf_splitterN113ton241n415_splitterN113ton414n415_9 , 0 , buf_splitterN113ton241n415_splitterN113ton414n415_8 );
buf_AQFP buf_splitterN113ton241n415_splitterN113ton414n415_7_( clk_5 , buf_splitterN113ton241n415_splitterN113ton414n415_8 , 0 , buf_splitterN113ton241n415_splitterN113ton414n415_7 );
buf_AQFP buf_splitterN113ton241n415_splitterN113ton414n415_6_( clk_7 , buf_splitterN113ton241n415_splitterN113ton414n415_7 , 0 , buf_splitterN113ton241n415_splitterN113ton414n415_6 );
buf_AQFP buf_splitterN113ton241n415_splitterN113ton414n415_5_( clk_1 , buf_splitterN113ton241n415_splitterN113ton414n415_6 , 0 , buf_splitterN113ton241n415_splitterN113ton414n415_5 );
buf_AQFP buf_splitterN113ton241n415_splitterN113ton414n415_4_( clk_3 , buf_splitterN113ton241n415_splitterN113ton414n415_5 , 0 , buf_splitterN113ton241n415_splitterN113ton414n415_4 );
buf_AQFP buf_splitterN113ton241n415_splitterN113ton414n415_3_( clk_5 , buf_splitterN113ton241n415_splitterN113ton414n415_4 , 0 , buf_splitterN113ton241n415_splitterN113ton414n415_3 );
buf_AQFP buf_splitterN113ton241n415_splitterN113ton414n415_2_( clk_7 , buf_splitterN113ton241n415_splitterN113ton414n415_3 , 0 , buf_splitterN113ton241n415_splitterN113ton414n415_2 );
buf_AQFP buf_splitterN113ton241n415_splitterN113ton414n415_1_( clk_1 , buf_splitterN113ton241n415_splitterN113ton414n415_2 , 0 , buf_splitterN113ton241n415_splitterN113ton414n415_1 );
buf_AQFP buf_splitterN117ton260n419_splitterN117ton418n419_10_( clk_7 , splitterN117ton260n419 , 0 , buf_splitterN117ton260n419_splitterN117ton418n419_10 );
buf_AQFP buf_splitterN117ton260n419_splitterN117ton418n419_9_( clk_1 , buf_splitterN117ton260n419_splitterN117ton418n419_10 , 0 , buf_splitterN117ton260n419_splitterN117ton418n419_9 );
buf_AQFP buf_splitterN117ton260n419_splitterN117ton418n419_8_( clk_3 , buf_splitterN117ton260n419_splitterN117ton418n419_9 , 0 , buf_splitterN117ton260n419_splitterN117ton418n419_8 );
buf_AQFP buf_splitterN117ton260n419_splitterN117ton418n419_7_( clk_5 , buf_splitterN117ton260n419_splitterN117ton418n419_8 , 0 , buf_splitterN117ton260n419_splitterN117ton418n419_7 );
buf_AQFP buf_splitterN117ton260n419_splitterN117ton418n419_6_( clk_7 , buf_splitterN117ton260n419_splitterN117ton418n419_7 , 0 , buf_splitterN117ton260n419_splitterN117ton418n419_6 );
buf_AQFP buf_splitterN117ton260n419_splitterN117ton418n419_5_( clk_1 , buf_splitterN117ton260n419_splitterN117ton418n419_6 , 0 , buf_splitterN117ton260n419_splitterN117ton418n419_5 );
buf_AQFP buf_splitterN117ton260n419_splitterN117ton418n419_4_( clk_3 , buf_splitterN117ton260n419_splitterN117ton418n419_5 , 0 , buf_splitterN117ton260n419_splitterN117ton418n419_4 );
buf_AQFP buf_splitterN117ton260n419_splitterN117ton418n419_3_( clk_5 , buf_splitterN117ton260n419_splitterN117ton418n419_4 , 0 , buf_splitterN117ton260n419_splitterN117ton418n419_3 );
buf_AQFP buf_splitterN117ton260n419_splitterN117ton418n419_2_( clk_7 , buf_splitterN117ton260n419_splitterN117ton418n419_3 , 0 , buf_splitterN117ton260n419_splitterN117ton418n419_2 );
buf_AQFP buf_splitterN117ton260n419_splitterN117ton418n419_1_( clk_1 , buf_splitterN117ton260n419_splitterN117ton418n419_2 , 0 , buf_splitterN117ton260n419_splitterN117ton418n419_1 );
buf_AQFP buf_splitterN121ton196n423_splitterN121ton422n423_11_( clk_5 , splitterN121ton196n423 , 0 , buf_splitterN121ton196n423_splitterN121ton422n423_11 );
buf_AQFP buf_splitterN121ton196n423_splitterN121ton422n423_10_( clk_7 , buf_splitterN121ton196n423_splitterN121ton422n423_11 , 0 , buf_splitterN121ton196n423_splitterN121ton422n423_10 );
buf_AQFP buf_splitterN121ton196n423_splitterN121ton422n423_9_( clk_1 , buf_splitterN121ton196n423_splitterN121ton422n423_10 , 0 , buf_splitterN121ton196n423_splitterN121ton422n423_9 );
buf_AQFP buf_splitterN121ton196n423_splitterN121ton422n423_8_( clk_3 , buf_splitterN121ton196n423_splitterN121ton422n423_9 , 0 , buf_splitterN121ton196n423_splitterN121ton422n423_8 );
buf_AQFP buf_splitterN121ton196n423_splitterN121ton422n423_7_( clk_5 , buf_splitterN121ton196n423_splitterN121ton422n423_8 , 0 , buf_splitterN121ton196n423_splitterN121ton422n423_7 );
buf_AQFP buf_splitterN121ton196n423_splitterN121ton422n423_6_( clk_7 , buf_splitterN121ton196n423_splitterN121ton422n423_7 , 0 , buf_splitterN121ton196n423_splitterN121ton422n423_6 );
buf_AQFP buf_splitterN121ton196n423_splitterN121ton422n423_5_( clk_1 , buf_splitterN121ton196n423_splitterN121ton422n423_6 , 0 , buf_splitterN121ton196n423_splitterN121ton422n423_5 );
buf_AQFP buf_splitterN121ton196n423_splitterN121ton422n423_4_( clk_3 , buf_splitterN121ton196n423_splitterN121ton422n423_5 , 0 , buf_splitterN121ton196n423_splitterN121ton422n423_4 );
buf_AQFP buf_splitterN121ton196n423_splitterN121ton422n423_3_( clk_5 , buf_splitterN121ton196n423_splitterN121ton422n423_4 , 0 , buf_splitterN121ton196n423_splitterN121ton422n423_3 );
buf_AQFP buf_splitterN121ton196n423_splitterN121ton422n423_2_( clk_7 , buf_splitterN121ton196n423_splitterN121ton422n423_3 , 0 , buf_splitterN121ton196n423_splitterN121ton422n423_2 );
buf_AQFP buf_splitterN121ton196n423_splitterN121ton422n423_1_( clk_1 , buf_splitterN121ton196n423_splitterN121ton422n423_2 , 0 , buf_splitterN121ton196n423_splitterN121ton422n423_1 );
buf_AQFP buf_splitterN125ton196n427_splitterN125ton426n427_11_( clk_5 , splitterN125ton196n427 , 0 , buf_splitterN125ton196n427_splitterN125ton426n427_11 );
buf_AQFP buf_splitterN125ton196n427_splitterN125ton426n427_10_( clk_7 , buf_splitterN125ton196n427_splitterN125ton426n427_11 , 0 , buf_splitterN125ton196n427_splitterN125ton426n427_10 );
buf_AQFP buf_splitterN125ton196n427_splitterN125ton426n427_9_( clk_1 , buf_splitterN125ton196n427_splitterN125ton426n427_10 , 0 , buf_splitterN125ton196n427_splitterN125ton426n427_9 );
buf_AQFP buf_splitterN125ton196n427_splitterN125ton426n427_8_( clk_3 , buf_splitterN125ton196n427_splitterN125ton426n427_9 , 0 , buf_splitterN125ton196n427_splitterN125ton426n427_8 );
buf_AQFP buf_splitterN125ton196n427_splitterN125ton426n427_7_( clk_5 , buf_splitterN125ton196n427_splitterN125ton426n427_8 , 0 , buf_splitterN125ton196n427_splitterN125ton426n427_7 );
buf_AQFP buf_splitterN125ton196n427_splitterN125ton426n427_6_( clk_7 , buf_splitterN125ton196n427_splitterN125ton426n427_7 , 0 , buf_splitterN125ton196n427_splitterN125ton426n427_6 );
buf_AQFP buf_splitterN125ton196n427_splitterN125ton426n427_5_( clk_1 , buf_splitterN125ton196n427_splitterN125ton426n427_6 , 0 , buf_splitterN125ton196n427_splitterN125ton426n427_5 );
buf_AQFP buf_splitterN125ton196n427_splitterN125ton426n427_4_( clk_3 , buf_splitterN125ton196n427_splitterN125ton426n427_5 , 0 , buf_splitterN125ton196n427_splitterN125ton426n427_4 );
buf_AQFP buf_splitterN125ton196n427_splitterN125ton426n427_3_( clk_5 , buf_splitterN125ton196n427_splitterN125ton426n427_4 , 0 , buf_splitterN125ton196n427_splitterN125ton426n427_3 );
buf_AQFP buf_splitterN125ton196n427_splitterN125ton426n427_2_( clk_7 , buf_splitterN125ton196n427_splitterN125ton426n427_3 , 0 , buf_splitterN125ton196n427_splitterN125ton426n427_2 );
buf_AQFP buf_splitterN125ton196n427_splitterN125ton426n427_1_( clk_1 , buf_splitterN125ton196n427_splitterN125ton426n427_2 , 0 , buf_splitterN125ton196n427_splitterN125ton426n427_1 );
buf_AQFP buf_splitterN13ton219n296_splitterN13ton295n296_11_( clk_7 , splitterN13ton219n296 , 0 , buf_splitterN13ton219n296_splitterN13ton295n296_11 );
buf_AQFP buf_splitterN13ton219n296_splitterN13ton295n296_10_( clk_1 , buf_splitterN13ton219n296_splitterN13ton295n296_11 , 0 , buf_splitterN13ton219n296_splitterN13ton295n296_10 );
buf_AQFP buf_splitterN13ton219n296_splitterN13ton295n296_9_( clk_3 , buf_splitterN13ton219n296_splitterN13ton295n296_10 , 0 , buf_splitterN13ton219n296_splitterN13ton295n296_9 );
buf_AQFP buf_splitterN13ton219n296_splitterN13ton295n296_8_( clk_5 , buf_splitterN13ton219n296_splitterN13ton295n296_9 , 0 , buf_splitterN13ton219n296_splitterN13ton295n296_8 );
buf_AQFP buf_splitterN13ton219n296_splitterN13ton295n296_7_( clk_7 , buf_splitterN13ton219n296_splitterN13ton295n296_8 , 0 , buf_splitterN13ton219n296_splitterN13ton295n296_7 );
buf_AQFP buf_splitterN13ton219n296_splitterN13ton295n296_6_( clk_1 , buf_splitterN13ton219n296_splitterN13ton295n296_7 , 0 , buf_splitterN13ton219n296_splitterN13ton295n296_6 );
buf_AQFP buf_splitterN13ton219n296_splitterN13ton295n296_5_( clk_3 , buf_splitterN13ton219n296_splitterN13ton295n296_6 , 0 , buf_splitterN13ton219n296_splitterN13ton295n296_5 );
buf_AQFP buf_splitterN13ton219n296_splitterN13ton295n296_4_( clk_5 , buf_splitterN13ton219n296_splitterN13ton295n296_5 , 0 , buf_splitterN13ton219n296_splitterN13ton295n296_4 );
buf_AQFP buf_splitterN13ton219n296_splitterN13ton295n296_3_( clk_7 , buf_splitterN13ton219n296_splitterN13ton295n296_4 , 0 , buf_splitterN13ton219n296_splitterN13ton295n296_3 );
buf_AQFP buf_splitterN13ton219n296_splitterN13ton295n296_2_( clk_1 , buf_splitterN13ton219n296_splitterN13ton295n296_3 , 0 , buf_splitterN13ton219n296_splitterN13ton295n296_2 );
buf_AQFP buf_splitterN13ton219n296_splitterN13ton295n296_1_( clk_3 , buf_splitterN13ton219n296_splitterN13ton295n296_2 , 0 , buf_splitterN13ton219n296_splitterN13ton295n296_1 );
buf_AQFP buf_splitterN17ton47n302_splitterN17ton301n302_12_( clk_5 , splitterN17ton47n302 , 0 , buf_splitterN17ton47n302_splitterN17ton301n302_12 );
buf_AQFP buf_splitterN17ton47n302_splitterN17ton301n302_11_( clk_7 , buf_splitterN17ton47n302_splitterN17ton301n302_12 , 0 , buf_splitterN17ton47n302_splitterN17ton301n302_11 );
buf_AQFP buf_splitterN17ton47n302_splitterN17ton301n302_10_( clk_1 , buf_splitterN17ton47n302_splitterN17ton301n302_11 , 0 , buf_splitterN17ton47n302_splitterN17ton301n302_10 );
buf_AQFP buf_splitterN17ton47n302_splitterN17ton301n302_9_( clk_3 , buf_splitterN17ton47n302_splitterN17ton301n302_10 , 0 , buf_splitterN17ton47n302_splitterN17ton301n302_9 );
buf_AQFP buf_splitterN17ton47n302_splitterN17ton301n302_8_( clk_5 , buf_splitterN17ton47n302_splitterN17ton301n302_9 , 0 , buf_splitterN17ton47n302_splitterN17ton301n302_8 );
buf_AQFP buf_splitterN17ton47n302_splitterN17ton301n302_7_( clk_7 , buf_splitterN17ton47n302_splitterN17ton301n302_8 , 0 , buf_splitterN17ton47n302_splitterN17ton301n302_7 );
buf_AQFP buf_splitterN17ton47n302_splitterN17ton301n302_6_( clk_1 , buf_splitterN17ton47n302_splitterN17ton301n302_7 , 0 , buf_splitterN17ton47n302_splitterN17ton301n302_6 );
buf_AQFP buf_splitterN17ton47n302_splitterN17ton301n302_5_( clk_3 , buf_splitterN17ton47n302_splitterN17ton301n302_6 , 0 , buf_splitterN17ton47n302_splitterN17ton301n302_5 );
buf_AQFP buf_splitterN17ton47n302_splitterN17ton301n302_4_( clk_5 , buf_splitterN17ton47n302_splitterN17ton301n302_5 , 0 , buf_splitterN17ton47n302_splitterN17ton301n302_4 );
buf_AQFP buf_splitterN17ton47n302_splitterN17ton301n302_3_( clk_7 , buf_splitterN17ton47n302_splitterN17ton301n302_4 , 0 , buf_splitterN17ton47n302_splitterN17ton301n302_3 );
buf_AQFP buf_splitterN17ton47n302_splitterN17ton301n302_2_( clk_1 , buf_splitterN17ton47n302_splitterN17ton301n302_3 , 0 , buf_splitterN17ton47n302_splitterN17ton301n302_2 );
buf_AQFP buf_splitterN17ton47n302_splitterN17ton301n302_1_( clk_3 , buf_splitterN17ton47n302_splitterN17ton301n302_2 , 0 , buf_splitterN17ton47n302_splitterN17ton301n302_1 );
buf_AQFP buf_splitterN21ton187n306_splitterN21ton305n306_12_( clk_5 , splitterN21ton187n306 , 0 , buf_splitterN21ton187n306_splitterN21ton305n306_12 );
buf_AQFP buf_splitterN21ton187n306_splitterN21ton305n306_11_( clk_7 , buf_splitterN21ton187n306_splitterN21ton305n306_12 , 0 , buf_splitterN21ton187n306_splitterN21ton305n306_11 );
buf_AQFP buf_splitterN21ton187n306_splitterN21ton305n306_10_( clk_1 , buf_splitterN21ton187n306_splitterN21ton305n306_11 , 0 , buf_splitterN21ton187n306_splitterN21ton305n306_10 );
buf_AQFP buf_splitterN21ton187n306_splitterN21ton305n306_9_( clk_3 , buf_splitterN21ton187n306_splitterN21ton305n306_10 , 0 , buf_splitterN21ton187n306_splitterN21ton305n306_9 );
buf_AQFP buf_splitterN21ton187n306_splitterN21ton305n306_8_( clk_5 , buf_splitterN21ton187n306_splitterN21ton305n306_9 , 0 , buf_splitterN21ton187n306_splitterN21ton305n306_8 );
buf_AQFP buf_splitterN21ton187n306_splitterN21ton305n306_7_( clk_7 , buf_splitterN21ton187n306_splitterN21ton305n306_8 , 0 , buf_splitterN21ton187n306_splitterN21ton305n306_7 );
buf_AQFP buf_splitterN21ton187n306_splitterN21ton305n306_6_( clk_1 , buf_splitterN21ton187n306_splitterN21ton305n306_7 , 0 , buf_splitterN21ton187n306_splitterN21ton305n306_6 );
buf_AQFP buf_splitterN21ton187n306_splitterN21ton305n306_5_( clk_3 , buf_splitterN21ton187n306_splitterN21ton305n306_6 , 0 , buf_splitterN21ton187n306_splitterN21ton305n306_5 );
buf_AQFP buf_splitterN21ton187n306_splitterN21ton305n306_4_( clk_5 , buf_splitterN21ton187n306_splitterN21ton305n306_5 , 0 , buf_splitterN21ton187n306_splitterN21ton305n306_4 );
buf_AQFP buf_splitterN21ton187n306_splitterN21ton305n306_3_( clk_7 , buf_splitterN21ton187n306_splitterN21ton305n306_4 , 0 , buf_splitterN21ton187n306_splitterN21ton305n306_3 );
buf_AQFP buf_splitterN21ton187n306_splitterN21ton305n306_2_( clk_1 , buf_splitterN21ton187n306_splitterN21ton305n306_3 , 0 , buf_splitterN21ton187n306_splitterN21ton305n306_2 );
buf_AQFP buf_splitterN21ton187n306_splitterN21ton305n306_1_( clk_3 , buf_splitterN21ton187n306_splitterN21ton305n306_2 , 0 , buf_splitterN21ton187n306_splitterN21ton305n306_1 );
buf_AQFP buf_splitterN25ton158n310_splitterN25ton309n310_11_( clk_7 , splitterN25ton158n310 , 0 , buf_splitterN25ton158n310_splitterN25ton309n310_11 );
buf_AQFP buf_splitterN25ton158n310_splitterN25ton309n310_10_( clk_1 , buf_splitterN25ton158n310_splitterN25ton309n310_11 , 0 , buf_splitterN25ton158n310_splitterN25ton309n310_10 );
buf_AQFP buf_splitterN25ton158n310_splitterN25ton309n310_9_( clk_3 , buf_splitterN25ton158n310_splitterN25ton309n310_10 , 0 , buf_splitterN25ton158n310_splitterN25ton309n310_9 );
buf_AQFP buf_splitterN25ton158n310_splitterN25ton309n310_8_( clk_5 , buf_splitterN25ton158n310_splitterN25ton309n310_9 , 0 , buf_splitterN25ton158n310_splitterN25ton309n310_8 );
buf_AQFP buf_splitterN25ton158n310_splitterN25ton309n310_7_( clk_7 , buf_splitterN25ton158n310_splitterN25ton309n310_8 , 0 , buf_splitterN25ton158n310_splitterN25ton309n310_7 );
buf_AQFP buf_splitterN25ton158n310_splitterN25ton309n310_6_( clk_1 , buf_splitterN25ton158n310_splitterN25ton309n310_7 , 0 , buf_splitterN25ton158n310_splitterN25ton309n310_6 );
buf_AQFP buf_splitterN25ton158n310_splitterN25ton309n310_5_( clk_3 , buf_splitterN25ton158n310_splitterN25ton309n310_6 , 0 , buf_splitterN25ton158n310_splitterN25ton309n310_5 );
buf_AQFP buf_splitterN25ton158n310_splitterN25ton309n310_4_( clk_5 , buf_splitterN25ton158n310_splitterN25ton309n310_5 , 0 , buf_splitterN25ton158n310_splitterN25ton309n310_4 );
buf_AQFP buf_splitterN25ton158n310_splitterN25ton309n310_3_( clk_7 , buf_splitterN25ton158n310_splitterN25ton309n310_4 , 0 , buf_splitterN25ton158n310_splitterN25ton309n310_3 );
buf_AQFP buf_splitterN25ton158n310_splitterN25ton309n310_2_( clk_1 , buf_splitterN25ton158n310_splitterN25ton309n310_3 , 0 , buf_splitterN25ton158n310_splitterN25ton309n310_2 );
buf_AQFP buf_splitterN25ton158n310_splitterN25ton309n310_1_( clk_3 , buf_splitterN25ton158n310_splitterN25ton309n310_2 , 0 , buf_splitterN25ton158n310_splitterN25ton309n310_1 );
buf_AQFP buf_splitterN29ton219n314_splitterN29ton313n314_11_( clk_7 , splitterN29ton219n314 , 0 , buf_splitterN29ton219n314_splitterN29ton313n314_11 );
buf_AQFP buf_splitterN29ton219n314_splitterN29ton313n314_10_( clk_1 , buf_splitterN29ton219n314_splitterN29ton313n314_11 , 0 , buf_splitterN29ton219n314_splitterN29ton313n314_10 );
buf_AQFP buf_splitterN29ton219n314_splitterN29ton313n314_9_( clk_3 , buf_splitterN29ton219n314_splitterN29ton313n314_10 , 0 , buf_splitterN29ton219n314_splitterN29ton313n314_9 );
buf_AQFP buf_splitterN29ton219n314_splitterN29ton313n314_8_( clk_5 , buf_splitterN29ton219n314_splitterN29ton313n314_9 , 0 , buf_splitterN29ton219n314_splitterN29ton313n314_8 );
buf_AQFP buf_splitterN29ton219n314_splitterN29ton313n314_7_( clk_7 , buf_splitterN29ton219n314_splitterN29ton313n314_8 , 0 , buf_splitterN29ton219n314_splitterN29ton313n314_7 );
buf_AQFP buf_splitterN29ton219n314_splitterN29ton313n314_6_( clk_1 , buf_splitterN29ton219n314_splitterN29ton313n314_7 , 0 , buf_splitterN29ton219n314_splitterN29ton313n314_6 );
buf_AQFP buf_splitterN29ton219n314_splitterN29ton313n314_5_( clk_3 , buf_splitterN29ton219n314_splitterN29ton313n314_6 , 0 , buf_splitterN29ton219n314_splitterN29ton313n314_5 );
buf_AQFP buf_splitterN29ton219n314_splitterN29ton313n314_4_( clk_5 , buf_splitterN29ton219n314_splitterN29ton313n314_5 , 0 , buf_splitterN29ton219n314_splitterN29ton313n314_4 );
buf_AQFP buf_splitterN29ton219n314_splitterN29ton313n314_3_( clk_7 , buf_splitterN29ton219n314_splitterN29ton313n314_4 , 0 , buf_splitterN29ton219n314_splitterN29ton313n314_3 );
buf_AQFP buf_splitterN29ton219n314_splitterN29ton313n314_2_( clk_1 , buf_splitterN29ton219n314_splitterN29ton313n314_3 , 0 , buf_splitterN29ton219n314_splitterN29ton313n314_2 );
buf_AQFP buf_splitterN29ton219n314_splitterN29ton313n314_1_( clk_3 , buf_splitterN29ton219n314_splitterN29ton313n314_2 , 0 , buf_splitterN29ton219n314_splitterN29ton313n314_1 );
buf_AQFP buf_splitterN33ton42n321_splitterN33ton320n321_11_( clk_7 , splitterN33ton42n321 , 0 , buf_splitterN33ton42n321_splitterN33ton320n321_11 );
buf_AQFP buf_splitterN33ton42n321_splitterN33ton320n321_10_( clk_1 , buf_splitterN33ton42n321_splitterN33ton320n321_11 , 0 , buf_splitterN33ton42n321_splitterN33ton320n321_10 );
buf_AQFP buf_splitterN33ton42n321_splitterN33ton320n321_9_( clk_3 , buf_splitterN33ton42n321_splitterN33ton320n321_10 , 0 , buf_splitterN33ton42n321_splitterN33ton320n321_9 );
buf_AQFP buf_splitterN33ton42n321_splitterN33ton320n321_8_( clk_5 , buf_splitterN33ton42n321_splitterN33ton320n321_9 , 0 , buf_splitterN33ton42n321_splitterN33ton320n321_8 );
buf_AQFP buf_splitterN33ton42n321_splitterN33ton320n321_7_( clk_7 , buf_splitterN33ton42n321_splitterN33ton320n321_8 , 0 , buf_splitterN33ton42n321_splitterN33ton320n321_7 );
buf_AQFP buf_splitterN33ton42n321_splitterN33ton320n321_6_( clk_1 , buf_splitterN33ton42n321_splitterN33ton320n321_7 , 0 , buf_splitterN33ton42n321_splitterN33ton320n321_6 );
buf_AQFP buf_splitterN33ton42n321_splitterN33ton320n321_5_( clk_3 , buf_splitterN33ton42n321_splitterN33ton320n321_6 , 0 , buf_splitterN33ton42n321_splitterN33ton320n321_5 );
buf_AQFP buf_splitterN33ton42n321_splitterN33ton320n321_4_( clk_5 , buf_splitterN33ton42n321_splitterN33ton320n321_5 , 0 , buf_splitterN33ton42n321_splitterN33ton320n321_4 );
buf_AQFP buf_splitterN33ton42n321_splitterN33ton320n321_3_( clk_7 , buf_splitterN33ton42n321_splitterN33ton320n321_4 , 0 , buf_splitterN33ton42n321_splitterN33ton320n321_3 );
buf_AQFP buf_splitterN33ton42n321_splitterN33ton320n321_2_( clk_1 , buf_splitterN33ton42n321_splitterN33ton320n321_3 , 0 , buf_splitterN33ton42n321_splitterN33ton320n321_2 );
buf_AQFP buf_splitterN33ton42n321_splitterN33ton320n321_1_( clk_3 , buf_splitterN33ton42n321_splitterN33ton320n321_2 , 0 , buf_splitterN33ton42n321_splitterN33ton320n321_1 );
buf_AQFP buf_splitterN37ton182n325_splitterN37ton324n325_11_( clk_7 , splitterN37ton182n325 , 0 , buf_splitterN37ton182n325_splitterN37ton324n325_11 );
buf_AQFP buf_splitterN37ton182n325_splitterN37ton324n325_10_( clk_1 , buf_splitterN37ton182n325_splitterN37ton324n325_11 , 0 , buf_splitterN37ton182n325_splitterN37ton324n325_10 );
buf_AQFP buf_splitterN37ton182n325_splitterN37ton324n325_9_( clk_3 , buf_splitterN37ton182n325_splitterN37ton324n325_10 , 0 , buf_splitterN37ton182n325_splitterN37ton324n325_9 );
buf_AQFP buf_splitterN37ton182n325_splitterN37ton324n325_8_( clk_5 , buf_splitterN37ton182n325_splitterN37ton324n325_9 , 0 , buf_splitterN37ton182n325_splitterN37ton324n325_8 );
buf_AQFP buf_splitterN37ton182n325_splitterN37ton324n325_7_( clk_7 , buf_splitterN37ton182n325_splitterN37ton324n325_8 , 0 , buf_splitterN37ton182n325_splitterN37ton324n325_7 );
buf_AQFP buf_splitterN37ton182n325_splitterN37ton324n325_6_( clk_1 , buf_splitterN37ton182n325_splitterN37ton324n325_7 , 0 , buf_splitterN37ton182n325_splitterN37ton324n325_6 );
buf_AQFP buf_splitterN37ton182n325_splitterN37ton324n325_5_( clk_3 , buf_splitterN37ton182n325_splitterN37ton324n325_6 , 0 , buf_splitterN37ton182n325_splitterN37ton324n325_5 );
buf_AQFP buf_splitterN37ton182n325_splitterN37ton324n325_4_( clk_5 , buf_splitterN37ton182n325_splitterN37ton324n325_5 , 0 , buf_splitterN37ton182n325_splitterN37ton324n325_4 );
buf_AQFP buf_splitterN37ton182n325_splitterN37ton324n325_3_( clk_7 , buf_splitterN37ton182n325_splitterN37ton324n325_4 , 0 , buf_splitterN37ton182n325_splitterN37ton324n325_3 );
buf_AQFP buf_splitterN37ton182n325_splitterN37ton324n325_2_( clk_1 , buf_splitterN37ton182n325_splitterN37ton324n325_3 , 0 , buf_splitterN37ton182n325_splitterN37ton324n325_2 );
buf_AQFP buf_splitterN37ton182n325_splitterN37ton324n325_1_( clk_3 , buf_splitterN37ton182n325_splitterN37ton324n325_2 , 0 , buf_splitterN37ton182n325_splitterN37ton324n325_1 );
buf_AQFP buf_splitterN41ton155n329_splitterN41ton328n329_11_( clk_7 , splitterN41ton155n329 , 0 , buf_splitterN41ton155n329_splitterN41ton328n329_11 );
buf_AQFP buf_splitterN41ton155n329_splitterN41ton328n329_10_( clk_1 , buf_splitterN41ton155n329_splitterN41ton328n329_11 , 0 , buf_splitterN41ton155n329_splitterN41ton328n329_10 );
buf_AQFP buf_splitterN41ton155n329_splitterN41ton328n329_9_( clk_3 , buf_splitterN41ton155n329_splitterN41ton328n329_10 , 0 , buf_splitterN41ton155n329_splitterN41ton328n329_9 );
buf_AQFP buf_splitterN41ton155n329_splitterN41ton328n329_8_( clk_5 , buf_splitterN41ton155n329_splitterN41ton328n329_9 , 0 , buf_splitterN41ton155n329_splitterN41ton328n329_8 );
buf_AQFP buf_splitterN41ton155n329_splitterN41ton328n329_7_( clk_7 , buf_splitterN41ton155n329_splitterN41ton328n329_8 , 0 , buf_splitterN41ton155n329_splitterN41ton328n329_7 );
buf_AQFP buf_splitterN41ton155n329_splitterN41ton328n329_6_( clk_1 , buf_splitterN41ton155n329_splitterN41ton328n329_7 , 0 , buf_splitterN41ton155n329_splitterN41ton328n329_6 );
buf_AQFP buf_splitterN41ton155n329_splitterN41ton328n329_5_( clk_3 , buf_splitterN41ton155n329_splitterN41ton328n329_6 , 0 , buf_splitterN41ton155n329_splitterN41ton328n329_5 );
buf_AQFP buf_splitterN41ton155n329_splitterN41ton328n329_4_( clk_5 , buf_splitterN41ton155n329_splitterN41ton328n329_5 , 0 , buf_splitterN41ton155n329_splitterN41ton328n329_4 );
buf_AQFP buf_splitterN41ton155n329_splitterN41ton328n329_3_( clk_7 , buf_splitterN41ton155n329_splitterN41ton328n329_4 , 0 , buf_splitterN41ton155n329_splitterN41ton328n329_3 );
buf_AQFP buf_splitterN41ton155n329_splitterN41ton328n329_2_( clk_1 , buf_splitterN41ton155n329_splitterN41ton328n329_3 , 0 , buf_splitterN41ton155n329_splitterN41ton328n329_2 );
buf_AQFP buf_splitterN41ton155n329_splitterN41ton328n329_1_( clk_3 , buf_splitterN41ton155n329_splitterN41ton328n329_2 , 0 , buf_splitterN41ton155n329_splitterN41ton328n329_1 );
buf_AQFP buf_splitterN45ton216n333_splitterN45ton332n333_11_( clk_7 , splitterN45ton216n333 , 0 , buf_splitterN45ton216n333_splitterN45ton332n333_11 );
buf_AQFP buf_splitterN45ton216n333_splitterN45ton332n333_10_( clk_1 , buf_splitterN45ton216n333_splitterN45ton332n333_11 , 0 , buf_splitterN45ton216n333_splitterN45ton332n333_10 );
buf_AQFP buf_splitterN45ton216n333_splitterN45ton332n333_9_( clk_3 , buf_splitterN45ton216n333_splitterN45ton332n333_10 , 0 , buf_splitterN45ton216n333_splitterN45ton332n333_9 );
buf_AQFP buf_splitterN45ton216n333_splitterN45ton332n333_8_( clk_5 , buf_splitterN45ton216n333_splitterN45ton332n333_9 , 0 , buf_splitterN45ton216n333_splitterN45ton332n333_8 );
buf_AQFP buf_splitterN45ton216n333_splitterN45ton332n333_7_( clk_7 , buf_splitterN45ton216n333_splitterN45ton332n333_8 , 0 , buf_splitterN45ton216n333_splitterN45ton332n333_7 );
buf_AQFP buf_splitterN45ton216n333_splitterN45ton332n333_6_( clk_1 , buf_splitterN45ton216n333_splitterN45ton332n333_7 , 0 , buf_splitterN45ton216n333_splitterN45ton332n333_6 );
buf_AQFP buf_splitterN45ton216n333_splitterN45ton332n333_5_( clk_3 , buf_splitterN45ton216n333_splitterN45ton332n333_6 , 0 , buf_splitterN45ton216n333_splitterN45ton332n333_5 );
buf_AQFP buf_splitterN45ton216n333_splitterN45ton332n333_4_( clk_5 , buf_splitterN45ton216n333_splitterN45ton332n333_5 , 0 , buf_splitterN45ton216n333_splitterN45ton332n333_4 );
buf_AQFP buf_splitterN45ton216n333_splitterN45ton332n333_3_( clk_7 , buf_splitterN45ton216n333_splitterN45ton332n333_4 , 0 , buf_splitterN45ton216n333_splitterN45ton332n333_3 );
buf_AQFP buf_splitterN45ton216n333_splitterN45ton332n333_2_( clk_1 , buf_splitterN45ton216n333_splitterN45ton332n333_3 , 0 , buf_splitterN45ton216n333_splitterN45ton332n333_2 );
buf_AQFP buf_splitterN45ton216n333_splitterN45ton332n333_1_( clk_3 , buf_splitterN45ton216n333_splitterN45ton332n333_2 , 0 , buf_splitterN45ton216n333_splitterN45ton332n333_1 );
buf_AQFP buf_splitterN49ton42n338_splitterN49ton337n338_11_( clk_7 , splitterN49ton42n338 , 0 , buf_splitterN49ton42n338_splitterN49ton337n338_11 );
buf_AQFP buf_splitterN49ton42n338_splitterN49ton337n338_10_( clk_1 , buf_splitterN49ton42n338_splitterN49ton337n338_11 , 0 , buf_splitterN49ton42n338_splitterN49ton337n338_10 );
buf_AQFP buf_splitterN49ton42n338_splitterN49ton337n338_9_( clk_3 , buf_splitterN49ton42n338_splitterN49ton337n338_10 , 0 , buf_splitterN49ton42n338_splitterN49ton337n338_9 );
buf_AQFP buf_splitterN49ton42n338_splitterN49ton337n338_8_( clk_5 , buf_splitterN49ton42n338_splitterN49ton337n338_9 , 0 , buf_splitterN49ton42n338_splitterN49ton337n338_8 );
buf_AQFP buf_splitterN49ton42n338_splitterN49ton337n338_7_( clk_7 , buf_splitterN49ton42n338_splitterN49ton337n338_8 , 0 , buf_splitterN49ton42n338_splitterN49ton337n338_7 );
buf_AQFP buf_splitterN49ton42n338_splitterN49ton337n338_6_( clk_1 , buf_splitterN49ton42n338_splitterN49ton337n338_7 , 0 , buf_splitterN49ton42n338_splitterN49ton337n338_6 );
buf_AQFP buf_splitterN49ton42n338_splitterN49ton337n338_5_( clk_3 , buf_splitterN49ton42n338_splitterN49ton337n338_6 , 0 , buf_splitterN49ton42n338_splitterN49ton337n338_5 );
buf_AQFP buf_splitterN49ton42n338_splitterN49ton337n338_4_( clk_5 , buf_splitterN49ton42n338_splitterN49ton337n338_5 , 0 , buf_splitterN49ton42n338_splitterN49ton337n338_4 );
buf_AQFP buf_splitterN49ton42n338_splitterN49ton337n338_3_( clk_7 , buf_splitterN49ton42n338_splitterN49ton337n338_4 , 0 , buf_splitterN49ton42n338_splitterN49ton337n338_3 );
buf_AQFP buf_splitterN49ton42n338_splitterN49ton337n338_2_( clk_1 , buf_splitterN49ton42n338_splitterN49ton337n338_3 , 0 , buf_splitterN49ton42n338_splitterN49ton337n338_2 );
buf_AQFP buf_splitterN49ton42n338_splitterN49ton337n338_1_( clk_3 , buf_splitterN49ton42n338_splitterN49ton337n338_2 , 0 , buf_splitterN49ton42n338_splitterN49ton337n338_1 );
buf_AQFP buf_splitterN5ton187n288_splitterN5ton287n288_12_( clk_5 , splitterN5ton187n288 , 0 , buf_splitterN5ton187n288_splitterN5ton287n288_12 );
buf_AQFP buf_splitterN5ton187n288_splitterN5ton287n288_11_( clk_7 , buf_splitterN5ton187n288_splitterN5ton287n288_12 , 0 , buf_splitterN5ton187n288_splitterN5ton287n288_11 );
buf_AQFP buf_splitterN5ton187n288_splitterN5ton287n288_10_( clk_1 , buf_splitterN5ton187n288_splitterN5ton287n288_11 , 0 , buf_splitterN5ton187n288_splitterN5ton287n288_10 );
buf_AQFP buf_splitterN5ton187n288_splitterN5ton287n288_9_( clk_3 , buf_splitterN5ton187n288_splitterN5ton287n288_10 , 0 , buf_splitterN5ton187n288_splitterN5ton287n288_9 );
buf_AQFP buf_splitterN5ton187n288_splitterN5ton287n288_8_( clk_5 , buf_splitterN5ton187n288_splitterN5ton287n288_9 , 0 , buf_splitterN5ton187n288_splitterN5ton287n288_8 );
buf_AQFP buf_splitterN5ton187n288_splitterN5ton287n288_7_( clk_7 , buf_splitterN5ton187n288_splitterN5ton287n288_8 , 0 , buf_splitterN5ton187n288_splitterN5ton287n288_7 );
buf_AQFP buf_splitterN5ton187n288_splitterN5ton287n288_6_( clk_1 , buf_splitterN5ton187n288_splitterN5ton287n288_7 , 0 , buf_splitterN5ton187n288_splitterN5ton287n288_6 );
buf_AQFP buf_splitterN5ton187n288_splitterN5ton287n288_5_( clk_3 , buf_splitterN5ton187n288_splitterN5ton287n288_6 , 0 , buf_splitterN5ton187n288_splitterN5ton287n288_5 );
buf_AQFP buf_splitterN5ton187n288_splitterN5ton287n288_4_( clk_5 , buf_splitterN5ton187n288_splitterN5ton287n288_5 , 0 , buf_splitterN5ton187n288_splitterN5ton287n288_4 );
buf_AQFP buf_splitterN5ton187n288_splitterN5ton287n288_3_( clk_7 , buf_splitterN5ton187n288_splitterN5ton287n288_4 , 0 , buf_splitterN5ton187n288_splitterN5ton287n288_3 );
buf_AQFP buf_splitterN5ton187n288_splitterN5ton287n288_2_( clk_1 , buf_splitterN5ton187n288_splitterN5ton287n288_3 , 0 , buf_splitterN5ton187n288_splitterN5ton287n288_2 );
buf_AQFP buf_splitterN5ton187n288_splitterN5ton287n288_1_( clk_3 , buf_splitterN5ton187n288_splitterN5ton287n288_2 , 0 , buf_splitterN5ton187n288_splitterN5ton287n288_1 );
buf_AQFP buf_splitterN53ton182n342_splitterN53ton341n342_11_( clk_7 , splitterN53ton182n342 , 0 , buf_splitterN53ton182n342_splitterN53ton341n342_11 );
buf_AQFP buf_splitterN53ton182n342_splitterN53ton341n342_10_( clk_1 , buf_splitterN53ton182n342_splitterN53ton341n342_11 , 0 , buf_splitterN53ton182n342_splitterN53ton341n342_10 );
buf_AQFP buf_splitterN53ton182n342_splitterN53ton341n342_9_( clk_3 , buf_splitterN53ton182n342_splitterN53ton341n342_10 , 0 , buf_splitterN53ton182n342_splitterN53ton341n342_9 );
buf_AQFP buf_splitterN53ton182n342_splitterN53ton341n342_8_( clk_5 , buf_splitterN53ton182n342_splitterN53ton341n342_9 , 0 , buf_splitterN53ton182n342_splitterN53ton341n342_8 );
buf_AQFP buf_splitterN53ton182n342_splitterN53ton341n342_7_( clk_7 , buf_splitterN53ton182n342_splitterN53ton341n342_8 , 0 , buf_splitterN53ton182n342_splitterN53ton341n342_7 );
buf_AQFP buf_splitterN53ton182n342_splitterN53ton341n342_6_( clk_1 , buf_splitterN53ton182n342_splitterN53ton341n342_7 , 0 , buf_splitterN53ton182n342_splitterN53ton341n342_6 );
buf_AQFP buf_splitterN53ton182n342_splitterN53ton341n342_5_( clk_3 , buf_splitterN53ton182n342_splitterN53ton341n342_6 , 0 , buf_splitterN53ton182n342_splitterN53ton341n342_5 );
buf_AQFP buf_splitterN53ton182n342_splitterN53ton341n342_4_( clk_5 , buf_splitterN53ton182n342_splitterN53ton341n342_5 , 0 , buf_splitterN53ton182n342_splitterN53ton341n342_4 );
buf_AQFP buf_splitterN53ton182n342_splitterN53ton341n342_3_( clk_7 , buf_splitterN53ton182n342_splitterN53ton341n342_4 , 0 , buf_splitterN53ton182n342_splitterN53ton341n342_3 );
buf_AQFP buf_splitterN53ton182n342_splitterN53ton341n342_2_( clk_1 , buf_splitterN53ton182n342_splitterN53ton341n342_3 , 0 , buf_splitterN53ton182n342_splitterN53ton341n342_2 );
buf_AQFP buf_splitterN53ton182n342_splitterN53ton341n342_1_( clk_3 , buf_splitterN53ton182n342_splitterN53ton341n342_2 , 0 , buf_splitterN53ton182n342_splitterN53ton341n342_1 );
buf_AQFP buf_splitterN57ton155n346_splitterN57ton345n346_11_( clk_7 , splitterN57ton155n346 , 0 , buf_splitterN57ton155n346_splitterN57ton345n346_11 );
buf_AQFP buf_splitterN57ton155n346_splitterN57ton345n346_10_( clk_1 , buf_splitterN57ton155n346_splitterN57ton345n346_11 , 0 , buf_splitterN57ton155n346_splitterN57ton345n346_10 );
buf_AQFP buf_splitterN57ton155n346_splitterN57ton345n346_9_( clk_3 , buf_splitterN57ton155n346_splitterN57ton345n346_10 , 0 , buf_splitterN57ton155n346_splitterN57ton345n346_9 );
buf_AQFP buf_splitterN57ton155n346_splitterN57ton345n346_8_( clk_5 , buf_splitterN57ton155n346_splitterN57ton345n346_9 , 0 , buf_splitterN57ton155n346_splitterN57ton345n346_8 );
buf_AQFP buf_splitterN57ton155n346_splitterN57ton345n346_7_( clk_7 , buf_splitterN57ton155n346_splitterN57ton345n346_8 , 0 , buf_splitterN57ton155n346_splitterN57ton345n346_7 );
buf_AQFP buf_splitterN57ton155n346_splitterN57ton345n346_6_( clk_1 , buf_splitterN57ton155n346_splitterN57ton345n346_7 , 0 , buf_splitterN57ton155n346_splitterN57ton345n346_6 );
buf_AQFP buf_splitterN57ton155n346_splitterN57ton345n346_5_( clk_3 , buf_splitterN57ton155n346_splitterN57ton345n346_6 , 0 , buf_splitterN57ton155n346_splitterN57ton345n346_5 );
buf_AQFP buf_splitterN57ton155n346_splitterN57ton345n346_4_( clk_5 , buf_splitterN57ton155n346_splitterN57ton345n346_5 , 0 , buf_splitterN57ton155n346_splitterN57ton345n346_4 );
buf_AQFP buf_splitterN57ton155n346_splitterN57ton345n346_3_( clk_7 , buf_splitterN57ton155n346_splitterN57ton345n346_4 , 0 , buf_splitterN57ton155n346_splitterN57ton345n346_3 );
buf_AQFP buf_splitterN57ton155n346_splitterN57ton345n346_2_( clk_1 , buf_splitterN57ton155n346_splitterN57ton345n346_3 , 0 , buf_splitterN57ton155n346_splitterN57ton345n346_2 );
buf_AQFP buf_splitterN57ton155n346_splitterN57ton345n346_1_( clk_3 , buf_splitterN57ton155n346_splitterN57ton345n346_2 , 0 , buf_splitterN57ton155n346_splitterN57ton345n346_1 );
buf_AQFP buf_splitterN61ton216n350_splitterN61ton349n350_11_( clk_7 , splitterN61ton216n350 , 0 , buf_splitterN61ton216n350_splitterN61ton349n350_11 );
buf_AQFP buf_splitterN61ton216n350_splitterN61ton349n350_10_( clk_1 , buf_splitterN61ton216n350_splitterN61ton349n350_11 , 0 , buf_splitterN61ton216n350_splitterN61ton349n350_10 );
buf_AQFP buf_splitterN61ton216n350_splitterN61ton349n350_9_( clk_3 , buf_splitterN61ton216n350_splitterN61ton349n350_10 , 0 , buf_splitterN61ton216n350_splitterN61ton349n350_9 );
buf_AQFP buf_splitterN61ton216n350_splitterN61ton349n350_8_( clk_5 , buf_splitterN61ton216n350_splitterN61ton349n350_9 , 0 , buf_splitterN61ton216n350_splitterN61ton349n350_8 );
buf_AQFP buf_splitterN61ton216n350_splitterN61ton349n350_7_( clk_7 , buf_splitterN61ton216n350_splitterN61ton349n350_8 , 0 , buf_splitterN61ton216n350_splitterN61ton349n350_7 );
buf_AQFP buf_splitterN61ton216n350_splitterN61ton349n350_6_( clk_1 , buf_splitterN61ton216n350_splitterN61ton349n350_7 , 0 , buf_splitterN61ton216n350_splitterN61ton349n350_6 );
buf_AQFP buf_splitterN61ton216n350_splitterN61ton349n350_5_( clk_3 , buf_splitterN61ton216n350_splitterN61ton349n350_6 , 0 , buf_splitterN61ton216n350_splitterN61ton349n350_5 );
buf_AQFP buf_splitterN61ton216n350_splitterN61ton349n350_4_( clk_5 , buf_splitterN61ton216n350_splitterN61ton349n350_5 , 0 , buf_splitterN61ton216n350_splitterN61ton349n350_4 );
buf_AQFP buf_splitterN61ton216n350_splitterN61ton349n350_3_( clk_7 , buf_splitterN61ton216n350_splitterN61ton349n350_4 , 0 , buf_splitterN61ton216n350_splitterN61ton349n350_3 );
buf_AQFP buf_splitterN61ton216n350_splitterN61ton349n350_2_( clk_1 , buf_splitterN61ton216n350_splitterN61ton349n350_3 , 0 , buf_splitterN61ton216n350_splitterN61ton349n350_2 );
buf_AQFP buf_splitterN61ton216n350_splitterN61ton349n350_1_( clk_3 , buf_splitterN61ton216n350_splitterN61ton349n350_2 , 0 , buf_splitterN61ton216n350_splitterN61ton349n350_1 );
buf_AQFP buf_splitterN65ton59n363_splitterN65ton362n363_11_( clk_5 , splitterN65ton59n363 , 0 , buf_splitterN65ton59n363_splitterN65ton362n363_11 );
buf_AQFP buf_splitterN65ton59n363_splitterN65ton362n363_10_( clk_7 , buf_splitterN65ton59n363_splitterN65ton362n363_11 , 0 , buf_splitterN65ton59n363_splitterN65ton362n363_10 );
buf_AQFP buf_splitterN65ton59n363_splitterN65ton362n363_9_( clk_1 , buf_splitterN65ton59n363_splitterN65ton362n363_10 , 0 , buf_splitterN65ton59n363_splitterN65ton362n363_9 );
buf_AQFP buf_splitterN65ton59n363_splitterN65ton362n363_8_( clk_3 , buf_splitterN65ton59n363_splitterN65ton362n363_9 , 0 , buf_splitterN65ton59n363_splitterN65ton362n363_8 );
buf_AQFP buf_splitterN65ton59n363_splitterN65ton362n363_7_( clk_5 , buf_splitterN65ton59n363_splitterN65ton362n363_8 , 0 , buf_splitterN65ton59n363_splitterN65ton362n363_7 );
buf_AQFP buf_splitterN65ton59n363_splitterN65ton362n363_6_( clk_7 , buf_splitterN65ton59n363_splitterN65ton362n363_7 , 0 , buf_splitterN65ton59n363_splitterN65ton362n363_6 );
buf_AQFP buf_splitterN65ton59n363_splitterN65ton362n363_5_( clk_1 , buf_splitterN65ton59n363_splitterN65ton362n363_6 , 0 , buf_splitterN65ton59n363_splitterN65ton362n363_5 );
buf_AQFP buf_splitterN65ton59n363_splitterN65ton362n363_4_( clk_3 , buf_splitterN65ton59n363_splitterN65ton362n363_5 , 0 , buf_splitterN65ton59n363_splitterN65ton362n363_4 );
buf_AQFP buf_splitterN65ton59n363_splitterN65ton362n363_3_( clk_5 , buf_splitterN65ton59n363_splitterN65ton362n363_4 , 0 , buf_splitterN65ton59n363_splitterN65ton362n363_3 );
buf_AQFP buf_splitterN65ton59n363_splitterN65ton362n363_2_( clk_7 , buf_splitterN65ton59n363_splitterN65ton362n363_3 , 0 , buf_splitterN65ton59n363_splitterN65ton362n363_2 );
buf_AQFP buf_splitterN65ton59n363_splitterN65ton362n363_1_( clk_1 , buf_splitterN65ton59n363_splitterN65ton362n363_2 , 0 , buf_splitterN65ton59n363_splitterN65ton362n363_1 );
buf_AQFP buf_splitterN69ton59n367_splitterN69ton366n367_11_( clk_5 , splitterN69ton59n367 , 0 , buf_splitterN69ton59n367_splitterN69ton366n367_11 );
buf_AQFP buf_splitterN69ton59n367_splitterN69ton366n367_10_( clk_7 , buf_splitterN69ton59n367_splitterN69ton366n367_11 , 0 , buf_splitterN69ton59n367_splitterN69ton366n367_10 );
buf_AQFP buf_splitterN69ton59n367_splitterN69ton366n367_9_( clk_1 , buf_splitterN69ton59n367_splitterN69ton366n367_10 , 0 , buf_splitterN69ton59n367_splitterN69ton366n367_9 );
buf_AQFP buf_splitterN69ton59n367_splitterN69ton366n367_8_( clk_3 , buf_splitterN69ton59n367_splitterN69ton366n367_9 , 0 , buf_splitterN69ton59n367_splitterN69ton366n367_8 );
buf_AQFP buf_splitterN69ton59n367_splitterN69ton366n367_7_( clk_5 , buf_splitterN69ton59n367_splitterN69ton366n367_8 , 0 , buf_splitterN69ton59n367_splitterN69ton366n367_7 );
buf_AQFP buf_splitterN69ton59n367_splitterN69ton366n367_6_( clk_7 , buf_splitterN69ton59n367_splitterN69ton366n367_7 , 0 , buf_splitterN69ton59n367_splitterN69ton366n367_6 );
buf_AQFP buf_splitterN69ton59n367_splitterN69ton366n367_5_( clk_1 , buf_splitterN69ton59n367_splitterN69ton366n367_6 , 0 , buf_splitterN69ton59n367_splitterN69ton366n367_5 );
buf_AQFP buf_splitterN69ton59n367_splitterN69ton366n367_4_( clk_3 , buf_splitterN69ton59n367_splitterN69ton366n367_5 , 0 , buf_splitterN69ton59n367_splitterN69ton366n367_4 );
buf_AQFP buf_splitterN69ton59n367_splitterN69ton366n367_3_( clk_5 , buf_splitterN69ton59n367_splitterN69ton366n367_4 , 0 , buf_splitterN69ton59n367_splitterN69ton366n367_3 );
buf_AQFP buf_splitterN69ton59n367_splitterN69ton366n367_2_( clk_7 , buf_splitterN69ton59n367_splitterN69ton366n367_3 , 0 , buf_splitterN69ton59n367_splitterN69ton366n367_2 );
buf_AQFP buf_splitterN69ton59n367_splitterN69ton366n367_1_( clk_1 , buf_splitterN69ton59n367_splitterN69ton366n367_2 , 0 , buf_splitterN69ton59n367_splitterN69ton366n367_1 );
buf_AQFP buf_splitterN73ton56n371_splitterN73ton370n371_11_( clk_5 , splitterN73ton56n371 , 0 , buf_splitterN73ton56n371_splitterN73ton370n371_11 );
buf_AQFP buf_splitterN73ton56n371_splitterN73ton370n371_10_( clk_7 , buf_splitterN73ton56n371_splitterN73ton370n371_11 , 0 , buf_splitterN73ton56n371_splitterN73ton370n371_10 );
buf_AQFP buf_splitterN73ton56n371_splitterN73ton370n371_9_( clk_1 , buf_splitterN73ton56n371_splitterN73ton370n371_10 , 0 , buf_splitterN73ton56n371_splitterN73ton370n371_9 );
buf_AQFP buf_splitterN73ton56n371_splitterN73ton370n371_8_( clk_3 , buf_splitterN73ton56n371_splitterN73ton370n371_9 , 0 , buf_splitterN73ton56n371_splitterN73ton370n371_8 );
buf_AQFP buf_splitterN73ton56n371_splitterN73ton370n371_7_( clk_5 , buf_splitterN73ton56n371_splitterN73ton370n371_8 , 0 , buf_splitterN73ton56n371_splitterN73ton370n371_7 );
buf_AQFP buf_splitterN73ton56n371_splitterN73ton370n371_6_( clk_7 , buf_splitterN73ton56n371_splitterN73ton370n371_7 , 0 , buf_splitterN73ton56n371_splitterN73ton370n371_6 );
buf_AQFP buf_splitterN73ton56n371_splitterN73ton370n371_5_( clk_1 , buf_splitterN73ton56n371_splitterN73ton370n371_6 , 0 , buf_splitterN73ton56n371_splitterN73ton370n371_5 );
buf_AQFP buf_splitterN73ton56n371_splitterN73ton370n371_4_( clk_3 , buf_splitterN73ton56n371_splitterN73ton370n371_5 , 0 , buf_splitterN73ton56n371_splitterN73ton370n371_4 );
buf_AQFP buf_splitterN73ton56n371_splitterN73ton370n371_3_( clk_5 , buf_splitterN73ton56n371_splitterN73ton370n371_4 , 0 , buf_splitterN73ton56n371_splitterN73ton370n371_3 );
buf_AQFP buf_splitterN73ton56n371_splitterN73ton370n371_2_( clk_7 , buf_splitterN73ton56n371_splitterN73ton370n371_3 , 0 , buf_splitterN73ton56n371_splitterN73ton370n371_2 );
buf_AQFP buf_splitterN73ton56n371_splitterN73ton370n371_1_( clk_1 , buf_splitterN73ton56n371_splitterN73ton370n371_2 , 0 , buf_splitterN73ton56n371_splitterN73ton370n371_1 );
buf_AQFP buf_splitterN77ton56n375_splitterN77ton374n375_11_( clk_5 , splitterN77ton56n375 , 0 , buf_splitterN77ton56n375_splitterN77ton374n375_11 );
buf_AQFP buf_splitterN77ton56n375_splitterN77ton374n375_10_( clk_7 , buf_splitterN77ton56n375_splitterN77ton374n375_11 , 0 , buf_splitterN77ton56n375_splitterN77ton374n375_10 );
buf_AQFP buf_splitterN77ton56n375_splitterN77ton374n375_9_( clk_1 , buf_splitterN77ton56n375_splitterN77ton374n375_10 , 0 , buf_splitterN77ton56n375_splitterN77ton374n375_9 );
buf_AQFP buf_splitterN77ton56n375_splitterN77ton374n375_8_( clk_3 , buf_splitterN77ton56n375_splitterN77ton374n375_9 , 0 , buf_splitterN77ton56n375_splitterN77ton374n375_8 );
buf_AQFP buf_splitterN77ton56n375_splitterN77ton374n375_7_( clk_5 , buf_splitterN77ton56n375_splitterN77ton374n375_8 , 0 , buf_splitterN77ton56n375_splitterN77ton374n375_7 );
buf_AQFP buf_splitterN77ton56n375_splitterN77ton374n375_6_( clk_7 , buf_splitterN77ton56n375_splitterN77ton374n375_7 , 0 , buf_splitterN77ton56n375_splitterN77ton374n375_6 );
buf_AQFP buf_splitterN77ton56n375_splitterN77ton374n375_5_( clk_1 , buf_splitterN77ton56n375_splitterN77ton374n375_6 , 0 , buf_splitterN77ton56n375_splitterN77ton374n375_5 );
buf_AQFP buf_splitterN77ton56n375_splitterN77ton374n375_4_( clk_3 , buf_splitterN77ton56n375_splitterN77ton374n375_5 , 0 , buf_splitterN77ton56n375_splitterN77ton374n375_4 );
buf_AQFP buf_splitterN77ton56n375_splitterN77ton374n375_3_( clk_5 , buf_splitterN77ton56n375_splitterN77ton374n375_4 , 0 , buf_splitterN77ton56n375_splitterN77ton374n375_3 );
buf_AQFP buf_splitterN77ton56n375_splitterN77ton374n375_2_( clk_7 , buf_splitterN77ton56n375_splitterN77ton374n375_3 , 0 , buf_splitterN77ton56n375_splitterN77ton374n375_2 );
buf_AQFP buf_splitterN77ton56n375_splitterN77ton374n375_1_( clk_1 , buf_splitterN77ton56n375_splitterN77ton374n375_2 , 0 , buf_splitterN77ton56n375_splitterN77ton374n375_1 );
buf_AQFP buf_splitterN81ton68n381_splitterN81ton380n381_11_( clk_5 , splitterN81ton68n381 , 0 , buf_splitterN81ton68n381_splitterN81ton380n381_11 );
buf_AQFP buf_splitterN81ton68n381_splitterN81ton380n381_10_( clk_7 , buf_splitterN81ton68n381_splitterN81ton380n381_11 , 0 , buf_splitterN81ton68n381_splitterN81ton380n381_10 );
buf_AQFP buf_splitterN81ton68n381_splitterN81ton380n381_9_( clk_1 , buf_splitterN81ton68n381_splitterN81ton380n381_10 , 0 , buf_splitterN81ton68n381_splitterN81ton380n381_9 );
buf_AQFP buf_splitterN81ton68n381_splitterN81ton380n381_8_( clk_3 , buf_splitterN81ton68n381_splitterN81ton380n381_9 , 0 , buf_splitterN81ton68n381_splitterN81ton380n381_8 );
buf_AQFP buf_splitterN81ton68n381_splitterN81ton380n381_7_( clk_5 , buf_splitterN81ton68n381_splitterN81ton380n381_8 , 0 , buf_splitterN81ton68n381_splitterN81ton380n381_7 );
buf_AQFP buf_splitterN81ton68n381_splitterN81ton380n381_6_( clk_7 , buf_splitterN81ton68n381_splitterN81ton380n381_7 , 0 , buf_splitterN81ton68n381_splitterN81ton380n381_6 );
buf_AQFP buf_splitterN81ton68n381_splitterN81ton380n381_5_( clk_1 , buf_splitterN81ton68n381_splitterN81ton380n381_6 , 0 , buf_splitterN81ton68n381_splitterN81ton380n381_5 );
buf_AQFP buf_splitterN81ton68n381_splitterN81ton380n381_4_( clk_3 , buf_splitterN81ton68n381_splitterN81ton380n381_5 , 0 , buf_splitterN81ton68n381_splitterN81ton380n381_4 );
buf_AQFP buf_splitterN81ton68n381_splitterN81ton380n381_3_( clk_5 , buf_splitterN81ton68n381_splitterN81ton380n381_4 , 0 , buf_splitterN81ton68n381_splitterN81ton380n381_3 );
buf_AQFP buf_splitterN81ton68n381_splitterN81ton380n381_2_( clk_7 , buf_splitterN81ton68n381_splitterN81ton380n381_3 , 0 , buf_splitterN81ton68n381_splitterN81ton380n381_2 );
buf_AQFP buf_splitterN81ton68n381_splitterN81ton380n381_1_( clk_1 , buf_splitterN81ton68n381_splitterN81ton380n381_2 , 0 , buf_splitterN81ton68n381_splitterN81ton380n381_1 );
buf_AQFP buf_splitterN85ton68n385_splitterN85ton384n385_11_( clk_5 , splitterN85ton68n385 , 0 , buf_splitterN85ton68n385_splitterN85ton384n385_11 );
buf_AQFP buf_splitterN85ton68n385_splitterN85ton384n385_10_( clk_7 , buf_splitterN85ton68n385_splitterN85ton384n385_11 , 0 , buf_splitterN85ton68n385_splitterN85ton384n385_10 );
buf_AQFP buf_splitterN85ton68n385_splitterN85ton384n385_9_( clk_1 , buf_splitterN85ton68n385_splitterN85ton384n385_10 , 0 , buf_splitterN85ton68n385_splitterN85ton384n385_9 );
buf_AQFP buf_splitterN85ton68n385_splitterN85ton384n385_8_( clk_3 , buf_splitterN85ton68n385_splitterN85ton384n385_9 , 0 , buf_splitterN85ton68n385_splitterN85ton384n385_8 );
buf_AQFP buf_splitterN85ton68n385_splitterN85ton384n385_7_( clk_5 , buf_splitterN85ton68n385_splitterN85ton384n385_8 , 0 , buf_splitterN85ton68n385_splitterN85ton384n385_7 );
buf_AQFP buf_splitterN85ton68n385_splitterN85ton384n385_6_( clk_7 , buf_splitterN85ton68n385_splitterN85ton384n385_7 , 0 , buf_splitterN85ton68n385_splitterN85ton384n385_6 );
buf_AQFP buf_splitterN85ton68n385_splitterN85ton384n385_5_( clk_1 , buf_splitterN85ton68n385_splitterN85ton384n385_6 , 0 , buf_splitterN85ton68n385_splitterN85ton384n385_5 );
buf_AQFP buf_splitterN85ton68n385_splitterN85ton384n385_4_( clk_3 , buf_splitterN85ton68n385_splitterN85ton384n385_5 , 0 , buf_splitterN85ton68n385_splitterN85ton384n385_4 );
buf_AQFP buf_splitterN85ton68n385_splitterN85ton384n385_3_( clk_5 , buf_splitterN85ton68n385_splitterN85ton384n385_4 , 0 , buf_splitterN85ton68n385_splitterN85ton384n385_3 );
buf_AQFP buf_splitterN85ton68n385_splitterN85ton384n385_2_( clk_7 , buf_splitterN85ton68n385_splitterN85ton384n385_3 , 0 , buf_splitterN85ton68n385_splitterN85ton384n385_2 );
buf_AQFP buf_splitterN85ton68n385_splitterN85ton384n385_1_( clk_1 , buf_splitterN85ton68n385_splitterN85ton384n385_2 , 0 , buf_splitterN85ton68n385_splitterN85ton384n385_1 );
buf_AQFP buf_splitterN89ton65n389_splitterN89ton388n389_11_( clk_5 , splitterN89ton65n389 , 0 , buf_splitterN89ton65n389_splitterN89ton388n389_11 );
buf_AQFP buf_splitterN89ton65n389_splitterN89ton388n389_10_( clk_7 , buf_splitterN89ton65n389_splitterN89ton388n389_11 , 0 , buf_splitterN89ton65n389_splitterN89ton388n389_10 );
buf_AQFP buf_splitterN89ton65n389_splitterN89ton388n389_9_( clk_1 , buf_splitterN89ton65n389_splitterN89ton388n389_10 , 0 , buf_splitterN89ton65n389_splitterN89ton388n389_9 );
buf_AQFP buf_splitterN89ton65n389_splitterN89ton388n389_8_( clk_3 , buf_splitterN89ton65n389_splitterN89ton388n389_9 , 0 , buf_splitterN89ton65n389_splitterN89ton388n389_8 );
buf_AQFP buf_splitterN89ton65n389_splitterN89ton388n389_7_( clk_5 , buf_splitterN89ton65n389_splitterN89ton388n389_8 , 0 , buf_splitterN89ton65n389_splitterN89ton388n389_7 );
buf_AQFP buf_splitterN89ton65n389_splitterN89ton388n389_6_( clk_7 , buf_splitterN89ton65n389_splitterN89ton388n389_7 , 0 , buf_splitterN89ton65n389_splitterN89ton388n389_6 );
buf_AQFP buf_splitterN89ton65n389_splitterN89ton388n389_5_( clk_1 , buf_splitterN89ton65n389_splitterN89ton388n389_6 , 0 , buf_splitterN89ton65n389_splitterN89ton388n389_5 );
buf_AQFP buf_splitterN89ton65n389_splitterN89ton388n389_4_( clk_3 , buf_splitterN89ton65n389_splitterN89ton388n389_5 , 0 , buf_splitterN89ton65n389_splitterN89ton388n389_4 );
buf_AQFP buf_splitterN89ton65n389_splitterN89ton388n389_3_( clk_5 , buf_splitterN89ton65n389_splitterN89ton388n389_4 , 0 , buf_splitterN89ton65n389_splitterN89ton388n389_3 );
buf_AQFP buf_splitterN89ton65n389_splitterN89ton388n389_2_( clk_7 , buf_splitterN89ton65n389_splitterN89ton388n389_3 , 0 , buf_splitterN89ton65n389_splitterN89ton388n389_2 );
buf_AQFP buf_splitterN89ton65n389_splitterN89ton388n389_1_( clk_1 , buf_splitterN89ton65n389_splitterN89ton388n389_2 , 0 , buf_splitterN89ton65n389_splitterN89ton388n389_1 );
buf_AQFP buf_splitterN9ton158n292_splitterN9ton291n292_11_( clk_7 , splitterN9ton158n292 , 0 , buf_splitterN9ton158n292_splitterN9ton291n292_11 );
buf_AQFP buf_splitterN9ton158n292_splitterN9ton291n292_10_( clk_1 , buf_splitterN9ton158n292_splitterN9ton291n292_11 , 0 , buf_splitterN9ton158n292_splitterN9ton291n292_10 );
buf_AQFP buf_splitterN9ton158n292_splitterN9ton291n292_9_( clk_3 , buf_splitterN9ton158n292_splitterN9ton291n292_10 , 0 , buf_splitterN9ton158n292_splitterN9ton291n292_9 );
buf_AQFP buf_splitterN9ton158n292_splitterN9ton291n292_8_( clk_5 , buf_splitterN9ton158n292_splitterN9ton291n292_9 , 0 , buf_splitterN9ton158n292_splitterN9ton291n292_8 );
buf_AQFP buf_splitterN9ton158n292_splitterN9ton291n292_7_( clk_7 , buf_splitterN9ton158n292_splitterN9ton291n292_8 , 0 , buf_splitterN9ton158n292_splitterN9ton291n292_7 );
buf_AQFP buf_splitterN9ton158n292_splitterN9ton291n292_6_( clk_1 , buf_splitterN9ton158n292_splitterN9ton291n292_7 , 0 , buf_splitterN9ton158n292_splitterN9ton291n292_6 );
buf_AQFP buf_splitterN9ton158n292_splitterN9ton291n292_5_( clk_3 , buf_splitterN9ton158n292_splitterN9ton291n292_6 , 0 , buf_splitterN9ton158n292_splitterN9ton291n292_5 );
buf_AQFP buf_splitterN9ton158n292_splitterN9ton291n292_4_( clk_5 , buf_splitterN9ton158n292_splitterN9ton291n292_5 , 0 , buf_splitterN9ton158n292_splitterN9ton291n292_4 );
buf_AQFP buf_splitterN9ton158n292_splitterN9ton291n292_3_( clk_7 , buf_splitterN9ton158n292_splitterN9ton291n292_4 , 0 , buf_splitterN9ton158n292_splitterN9ton291n292_3 );
buf_AQFP buf_splitterN9ton158n292_splitterN9ton291n292_2_( clk_1 , buf_splitterN9ton158n292_splitterN9ton291n292_3 , 0 , buf_splitterN9ton158n292_splitterN9ton291n292_2 );
buf_AQFP buf_splitterN9ton158n292_splitterN9ton291n292_1_( clk_3 , buf_splitterN9ton158n292_splitterN9ton291n292_2 , 0 , buf_splitterN9ton158n292_splitterN9ton291n292_1 );
buf_AQFP buf_splitterN93ton65n393_splitterN93ton392n393_11_( clk_5 , splitterN93ton65n393 , 0 , buf_splitterN93ton65n393_splitterN93ton392n393_11 );
buf_AQFP buf_splitterN93ton65n393_splitterN93ton392n393_10_( clk_7 , buf_splitterN93ton65n393_splitterN93ton392n393_11 , 0 , buf_splitterN93ton65n393_splitterN93ton392n393_10 );
buf_AQFP buf_splitterN93ton65n393_splitterN93ton392n393_9_( clk_1 , buf_splitterN93ton65n393_splitterN93ton392n393_10 , 0 , buf_splitterN93ton65n393_splitterN93ton392n393_9 );
buf_AQFP buf_splitterN93ton65n393_splitterN93ton392n393_8_( clk_3 , buf_splitterN93ton65n393_splitterN93ton392n393_9 , 0 , buf_splitterN93ton65n393_splitterN93ton392n393_8 );
buf_AQFP buf_splitterN93ton65n393_splitterN93ton392n393_7_( clk_5 , buf_splitterN93ton65n393_splitterN93ton392n393_8 , 0 , buf_splitterN93ton65n393_splitterN93ton392n393_7 );
buf_AQFP buf_splitterN93ton65n393_splitterN93ton392n393_6_( clk_7 , buf_splitterN93ton65n393_splitterN93ton392n393_7 , 0 , buf_splitterN93ton65n393_splitterN93ton392n393_6 );
buf_AQFP buf_splitterN93ton65n393_splitterN93ton392n393_5_( clk_1 , buf_splitterN93ton65n393_splitterN93ton392n393_6 , 0 , buf_splitterN93ton65n393_splitterN93ton392n393_5 );
buf_AQFP buf_splitterN93ton65n393_splitterN93ton392n393_4_( clk_3 , buf_splitterN93ton65n393_splitterN93ton392n393_5 , 0 , buf_splitterN93ton65n393_splitterN93ton392n393_4 );
buf_AQFP buf_splitterN93ton65n393_splitterN93ton392n393_3_( clk_5 , buf_splitterN93ton65n393_splitterN93ton392n393_4 , 0 , buf_splitterN93ton65n393_splitterN93ton392n393_3 );
buf_AQFP buf_splitterN93ton65n393_splitterN93ton392n393_2_( clk_7 , buf_splitterN93ton65n393_splitterN93ton392n393_3 , 0 , buf_splitterN93ton65n393_splitterN93ton392n393_2 );
buf_AQFP buf_splitterN93ton65n393_splitterN93ton392n393_1_( clk_1 , buf_splitterN93ton65n393_splitterN93ton392n393_2 , 0 , buf_splitterN93ton65n393_splitterN93ton392n393_1 );
buf_AQFP buf_splitterN97ton241n398_splitterN97ton397n398_10_( clk_7 , splitterN97ton241n398 , 0 , buf_splitterN97ton241n398_splitterN97ton397n398_10 );
buf_AQFP buf_splitterN97ton241n398_splitterN97ton397n398_9_( clk_1 , buf_splitterN97ton241n398_splitterN97ton397n398_10 , 0 , buf_splitterN97ton241n398_splitterN97ton397n398_9 );
buf_AQFP buf_splitterN97ton241n398_splitterN97ton397n398_8_( clk_3 , buf_splitterN97ton241n398_splitterN97ton397n398_9 , 0 , buf_splitterN97ton241n398_splitterN97ton397n398_8 );
buf_AQFP buf_splitterN97ton241n398_splitterN97ton397n398_7_( clk_5 , buf_splitterN97ton241n398_splitterN97ton397n398_8 , 0 , buf_splitterN97ton241n398_splitterN97ton397n398_7 );
buf_AQFP buf_splitterN97ton241n398_splitterN97ton397n398_6_( clk_7 , buf_splitterN97ton241n398_splitterN97ton397n398_7 , 0 , buf_splitterN97ton241n398_splitterN97ton397n398_6 );
buf_AQFP buf_splitterN97ton241n398_splitterN97ton397n398_5_( clk_1 , buf_splitterN97ton241n398_splitterN97ton397n398_6 , 0 , buf_splitterN97ton241n398_splitterN97ton397n398_5 );
buf_AQFP buf_splitterN97ton241n398_splitterN97ton397n398_4_( clk_3 , buf_splitterN97ton241n398_splitterN97ton397n398_5 , 0 , buf_splitterN97ton241n398_splitterN97ton397n398_4 );
buf_AQFP buf_splitterN97ton241n398_splitterN97ton397n398_3_( clk_5 , buf_splitterN97ton241n398_splitterN97ton397n398_4 , 0 , buf_splitterN97ton241n398_splitterN97ton397n398_3 );
buf_AQFP buf_splitterN97ton241n398_splitterN97ton397n398_2_( clk_7 , buf_splitterN97ton241n398_splitterN97ton397n398_3 , 0 , buf_splitterN97ton241n398_splitterN97ton397n398_2 );
buf_AQFP buf_splitterN97ton241n398_splitterN97ton397n398_1_( clk_1 , buf_splitterN97ton241n398_splitterN97ton397n398_2 , 0 , buf_splitterN97ton241n398_splitterN97ton397n398_1 );
buf_AQFP buf_splittern78ton238n336_splittern78ton282n336_4_( clk_3 , splittern78ton238n336 , 0 , buf_splittern78ton238n336_splittern78ton282n336_4 );
buf_AQFP buf_splittern78ton238n336_splittern78ton282n336_3_( clk_5 , buf_splittern78ton238n336_splittern78ton282n336_4 , 0 , buf_splittern78ton238n336_splittern78ton282n336_3 );
buf_AQFP buf_splittern78ton238n336_splittern78ton282n336_2_( clk_7 , buf_splittern78ton238n336_splittern78ton282n336_3 , 0 , buf_splittern78ton238n336_splittern78ton282n336_2 );
buf_AQFP buf_splittern78ton238n336_splittern78ton282n336_1_( clk_1 , buf_splittern78ton238n336_splittern78ton282n336_2 , 0 , buf_splittern78ton238n336_splittern78ton282n336_1 );
buf_AQFP buf_splittern115ton353n421_splittern115ton369n421_3_( clk_3 , splittern115ton353n421 , 0 , buf_splittern115ton353n421_splittern115ton369n421_3 );
buf_AQFP buf_splittern115ton353n421_splittern115ton369n421_2_( clk_5 , buf_splittern115ton353n421_splittern115ton369n421_3 , 0 , buf_splittern115ton353n421_splittern115ton369n421_2 );
buf_AQFP buf_splittern115ton353n421_splittern115ton369n421_1_( clk_7 , buf_splittern115ton353n421_splittern115ton369n421_2 , 0 , buf_splittern115ton353n421_splittern115ton369n421_1 );
buf_AQFP buf_splittern152ton353n425_splittern152ton373n425_3_( clk_3 , splittern152ton353n425 , 0 , buf_splittern152ton353n425_splittern152ton373n425_3 );
buf_AQFP buf_splittern152ton353n425_splittern152ton373n425_2_( clk_5 , buf_splittern152ton353n425_splittern152ton373n425_3 , 0 , buf_splittern152ton353n425_splittern152ton373n425_2 );
buf_AQFP buf_splittern152ton353n425_splittern152ton373n425_1_( clk_7 , buf_splittern152ton353n425_splittern152ton373n425_2 , 0 , buf_splittern152ton353n425_splittern152ton373n425_1 );
buf_AQFP buf_splittern153ton355n318_splittern153ton281n318_3_( clk_3 , splittern153ton355n318 , 0 , buf_splittern153ton355n318_splittern153ton281n318_3 );
buf_AQFP buf_splittern153ton355n318_splittern153ton281n318_2_( clk_5 , buf_splittern153ton355n318_splittern153ton281n318_3 , 0 , buf_splittern153ton355n318_splittern153ton281n318_2 );
buf_AQFP buf_splittern153ton355n318_splittern153ton281n318_1_( clk_7 , buf_splittern153ton355n318_splittern153ton281n318_2 , 0 , buf_splittern153ton355n318_splittern153ton281n318_1 );
buf_AQFP buf_splittern181ton236n344_splittern181ton290n344_3_( clk_4 , splittern181ton236n344 , 0 , buf_splittern181ton236n344_splittern181ton290n344_3 );
buf_AQFP buf_splittern181ton236n344_splittern181ton290n344_2_( clk_6 , buf_splittern181ton236n344_splittern181ton290n344_3 , 0 , buf_splittern181ton236n344_splittern181ton290n344_2 );
buf_AQFP buf_splittern181ton236n344_splittern181ton290n344_1_( clk_8 , buf_splittern181ton236n344_splittern181ton290n344_2 , 0 , buf_splittern181ton236n344_splittern181ton290n344_1 );
buf_AQFP buf_splittern209ton210n340_splittern209ton238n340_1_( clk_1 , splittern209ton210n340 , 0 , buf_splittern209ton210n340_splittern209ton238n340_1 );
buf_AQFP buf_splittern209ton238n340_splittern209ton286n340_3_( clk_4 , splittern209ton238n340 , 0 , buf_splittern209ton238n340_splittern209ton286n340_3 );
buf_AQFP buf_splittern209ton238n340_splittern209ton286n340_2_( clk_6 , buf_splittern209ton238n340_splittern209ton286n340_3 , 0 , buf_splittern209ton238n340_splittern209ton286n340_2 );
buf_AQFP buf_splittern209ton238n340_splittern209ton286n340_1_( clk_8 , buf_splittern209ton238n340_splittern209ton286n340_2 , 0 , buf_splittern209ton238n340_splittern209ton286n340_1 );
buf_AQFP buf_splitterfromn210_n395_3_( clk_3 , splitterfromn210 , 0 , buf_splitterfromn210_n395_3 );
buf_AQFP buf_splitterfromn210_n395_2_( clk_5 , buf_splitterfromn210_n395_3 , 0 , buf_splitterfromn210_n395_2 );
buf_AQFP buf_splitterfromn210_n395_1_( clk_7 , buf_splitterfromn210_n395_2 , 0 , buf_splitterfromn210_n395_1 );
buf_AQFP buf_splitterfromn211_n412_2_( clk_5 , splitterfromn211 , 0 , buf_splitterfromn211_n412_2 );
buf_AQFP buf_splitterfromn211_n412_1_( clk_7 , buf_splitterfromn211_n412_2 , 0 , buf_splitterfromn211_n412_1 );
buf_AQFP buf_splitterfromn212_n360_3_( clk_3 , splitterfromn212 , 0 , buf_splitterfromn212_n360_3 );
buf_AQFP buf_splitterfromn212_n360_2_( clk_5 , buf_splitterfromn212_n360_3 , 0 , buf_splitterfromn212_n360_2 );
buf_AQFP buf_splitterfromn212_n360_1_( clk_7 , buf_splitterfromn212_n360_2 , 0 , buf_splitterfromn212_n360_1 );
buf_AQFP buf_splitterfromn213_n378_2_( clk_5 , splitterfromn213 , 0 , buf_splitterfromn213_n378_2 );
buf_AQFP buf_splitterfromn213_n378_1_( clk_7 , buf_splitterfromn213_n378_2 , 0 , buf_splitterfromn213_n378_1 );
buf_AQFP buf_splittern233ton234n348_splittern233ton294n348_2_( clk_6 , splittern233ton234n348 , 0 , buf_splittern233ton234n348_splittern233ton294n348_2 );
buf_AQFP buf_splittern233ton234n348_splittern233ton294n348_1_( clk_8 , buf_splittern233ton234n348_splittern233ton294n348_2 , 0 , buf_splittern233ton234n348_splittern233ton294n348_1 );
buf_AQFP buf_splitterfromn235_n359_1_( clk_5 , splitterfromn235 , 0 , buf_splitterfromn235_n359_1 );
buf_AQFP buf_splittern259ton356n413_splittern259ton361n413_3_( clk_3 , splittern259ton356n413 , 0 , buf_splittern259ton356n413_splittern259ton361n413_3 );
buf_AQFP buf_splittern259ton356n413_splittern259ton361n413_2_( clk_5 , buf_splittern259ton356n413_splittern259ton361n413_3 , 0 , buf_splittern259ton356n413_splittern259ton361n413_2 );
buf_AQFP buf_splittern259ton356n413_splittern259ton361n413_1_( clk_7 , buf_splittern259ton356n413_splittern259ton361n413_2 , 0 , buf_splittern259ton356n413_splittern259ton361n413_1 );
buf_AQFP buf_splittern278ton356n417_splittern278ton365n417_3_( clk_3 , splittern278ton356n417 , 0 , buf_splittern278ton356n417_splittern278ton365n417_3 );
buf_AQFP buf_splittern278ton356n417_splittern278ton365n417_2_( clk_5 , buf_splittern278ton356n417_splittern278ton365n417_3 , 0 , buf_splittern278ton356n417_splittern278ton365n417_2 );
buf_AQFP buf_splittern278ton356n417_splittern278ton365n417_1_( clk_7 , buf_splittern278ton356n417_splittern278ton365n417_2 , 0 , buf_splittern278ton356n417_splittern278ton365n417_1 );
buf_AQFP buf_splitterfromn279_n280_3_( clk_3 , splitterfromn279 , 0 , buf_splitterfromn279_n280_3 );
buf_AQFP buf_splitterfromn279_n280_2_( clk_5 , buf_splitterfromn279_n280_3 , 0 , buf_splitterfromn279_n280_2 );
buf_AQFP buf_splitterfromn279_n280_1_( clk_7 , buf_splitterfromn279_n280_2 , 0 , buf_splitterfromn279_n280_1 );
buf_AQFP buf_splittern298ton355n335_splittern298ton299n335_3_( clk_3 , splittern298ton355n335 , 0 , buf_splittern298ton355n335_splittern298ton299n335_3 );
buf_AQFP buf_splittern298ton355n335_splittern298ton299n335_2_( clk_5 , buf_splittern298ton355n335_splittern298ton299n335_3 , 0 , buf_splittern298ton355n335_splittern298ton299n335_2 );
buf_AQFP buf_splittern298ton355n335_splittern298ton299n335_1_( clk_7 , buf_splittern298ton355n335_splittern298ton299n335_2 , 0 , buf_splittern298ton355n335_splittern298ton299n335_1 );
buf_AQFP buf_splitterfromn316_n317_3_( clk_3 , splitterfromn316 , 0 , buf_splitterfromn316_n317_3 );
buf_AQFP buf_splitterfromn316_n317_2_( clk_5 , buf_splitterfromn316_n317_3 , 0 , buf_splitterfromn316_n317_2 );
buf_AQFP buf_splitterfromn316_n317_1_( clk_7 , buf_splitterfromn316_n317_2 , 0 , buf_splitterfromn316_n317_1 );
splitter_AQFP splitterN1ton46n284_( clk_2 , N1 , 0 , splitterN1ton46n284 );
splitter_AQFP splitterN1ton47n284_( clk_3 , splitterN1ton46n284 , 0 , splitterN1ton47n284 );
splitter_AQFP splitterN1ton283n284_( clk_4 , buf_splitterN1ton47n284_splitterN1ton283n284_1 , 0 , splitterN1ton283n284 );
splitter_AQFP splitterN101ton170n402_( clk_3 , N101 , 0 , splitterN101ton170n402 );
splitter_AQFP splitterN101ton260n402_( clk_5 , splitterN101ton170n402 , 0 , splitterN101ton260n402 );
splitter_AQFP splitterN101ton401n402_( clk_2 , buf_splitterN101ton260n402_splitterN101ton401n402_1 , 0 , splitterN101ton401n402 );
splitter_AQFP splitterN105ton167n406_( clk_2 , N105 , 0 , splitterN105ton167n406 );
splitter_AQFP splitterN105ton168n406_( clk_3 , splitterN105ton167n406 , 0 , splitterN105ton168n406 );
splitter_AQFP splitterN105ton405n406_( clk_2 , buf_splitterN105ton168n406_splitterN105ton405n406_1 , 0 , splitterN105ton405n406 );
splitter_AQFP splitterN109ton117n410_( clk_2 , N109 , 0 , splitterN109ton117n410 );
splitter_AQFP splitterN109ton168n410_( clk_3 , splitterN109ton117n410 , 0 , splitterN109ton168n410 );
splitter_AQFP splitterN109ton409n410_( clk_2 , buf_splitterN109ton168n410_splitterN109ton409n410_1 , 0 , splitterN109ton409n410 );
splitter_AQFP splitterN113ton198n415_( clk_3 , N113 , 0 , splitterN113ton198n415 );
splitter_AQFP splitterN113ton241n415_( clk_5 , splitterN113ton198n415 , 0 , splitterN113ton241n415 );
splitter_AQFP splitterN113ton414n415_( clk_2 , buf_splitterN113ton241n415_splitterN113ton414n415_1 , 0 , splitterN113ton414n415 );
splitter_AQFP splitterN117ton198n419_( clk_3 , N117 , 0 , splitterN117ton198n419 );
splitter_AQFP splitterN117ton260n419_( clk_5 , splitterN117ton198n419 , 0 , splitterN117ton260n419 );
splitter_AQFP splitterN117ton418n419_( clk_2 , buf_splitterN117ton260n419_splitterN117ton418n419_1 , 0 , splitterN117ton418n419 );
splitter_AQFP splitterN121ton195n423_( clk_2 , N121 , 0 , splitterN121ton195n423 );
splitter_AQFP splitterN121ton196n423_( clk_3 , splitterN121ton195n423 , 0 , splitterN121ton196n423 );
splitter_AQFP splitterN121ton422n423_( clk_2 , buf_splitterN121ton196n423_splitterN121ton422n423_1 , 0 , splitterN121ton422n423 );
splitter_AQFP splitterN125ton117n427_( clk_2 , N125 , 0 , splitterN125ton117n427 );
splitter_AQFP splitterN125ton196n427_( clk_3 , splitterN125ton117n427 , 0 , splitterN125ton196n427 );
splitter_AQFP splitterN125ton426n427_( clk_2 , buf_splitterN125ton196n427_splitterN125ton426n427_1 , 0 , splitterN125ton426n427 );
splitter_AQFP splitterN13ton92n296_( clk_3 , N13 , 0 , splitterN13ton92n296 );
splitter_AQFP splitterN13ton219n296_( clk_5 , splitterN13ton92n296 , 0 , splitterN13ton219n296 );
splitter_AQFP splitterN13ton295n296_( clk_4 , buf_splitterN13ton219n296_splitterN13ton295n296_1 , 0 , splitterN13ton295n296 );
splitter_AQFP splitterN137ton116n79_( clk_2 , N137 , 0 , splitterN137ton116n79 );
splitter_AQFP splitterN137ton185n79_( clk_3 , splitterN137ton116n79 , 0 , splitterN137ton185n79 );
splitter_AQFP splitterN137ton154n79_( clk_4 , splitterN137ton185n79 , 0 , splitterN137ton154n79 );
splitter_AQFP splitterN17ton132n302_( clk_2 , N17 , 0 , splitterN17ton132n302 );
splitter_AQFP splitterN17ton47n302_( clk_3 , splitterN17ton132n302 , 0 , splitterN17ton47n302 );
splitter_AQFP splitterN17ton301n302_( clk_4 , buf_splitterN17ton47n302_splitterN17ton301n302_1 , 0 , splitterN17ton301n302 );
splitter_AQFP splitterN21ton132n306_( clk_2 , N21 , 0 , splitterN21ton132n306 );
splitter_AQFP splitterN21ton187n306_( clk_3 , splitterN21ton132n306 , 0 , splitterN21ton187n306 );
splitter_AQFP splitterN21ton305n306_( clk_4 , buf_splitterN21ton187n306_splitterN21ton305n306_1 , 0 , splitterN21ton305n306 );
splitter_AQFP splitterN25ton129n310_( clk_3 , N25 , 0 , splitterN25ton129n310 );
splitter_AQFP splitterN25ton158n310_( clk_5 , splitterN25ton129n310 , 0 , splitterN25ton158n310 );
splitter_AQFP splitterN25ton309n310_( clk_4 , buf_splitterN25ton158n310_splitterN25ton309n310_1 , 0 , splitterN25ton309n310 );
splitter_AQFP splitterN29ton129n314_( clk_3 , N29 , 0 , splitterN29ton129n314 );
splitter_AQFP splitterN29ton219n314_( clk_5 , splitterN29ton129n314 , 0 , splitterN29ton219n314 );
splitter_AQFP splitterN29ton313n314_( clk_4 , buf_splitterN29ton219n314_splitterN29ton313n314_1 , 0 , splitterN29ton313n314 );
splitter_AQFP splitterN33ton104n321_( clk_3 , N33 , 0 , splitterN33ton104n321 );
splitter_AQFP splitterN33ton42n321_( clk_5 , splitterN33ton104n321 , 0 , splitterN33ton42n321 );
splitter_AQFP splitterN33ton320n321_( clk_4 , buf_splitterN33ton42n321_splitterN33ton320n321_1 , 0 , splitterN33ton320n321 );
splitter_AQFP splitterN37ton104n325_( clk_3 , N37 , 0 , splitterN37ton104n325 );
splitter_AQFP splitterN37ton182n325_( clk_5 , splitterN37ton104n325 , 0 , splitterN37ton182n325 );
splitter_AQFP splitterN37ton324n325_( clk_4 , buf_splitterN37ton182n325_splitterN37ton324n325_1 , 0 , splitterN37ton324n325 );
splitter_AQFP splitterN41ton101n329_( clk_3 , N41 , 0 , splitterN41ton101n329 );
splitter_AQFP splitterN41ton155n329_( clk_5 , splitterN41ton101n329 , 0 , splitterN41ton155n329 );
splitter_AQFP splitterN41ton328n329_( clk_4 , buf_splitterN41ton155n329_splitterN41ton328n329_1 , 0 , splitterN41ton328n329 );
splitter_AQFP splitterN45ton101n333_( clk_3 , N45 , 0 , splitterN45ton101n333 );
splitter_AQFP splitterN45ton216n333_( clk_5 , splitterN45ton101n333 , 0 , splitterN45ton216n333 );
splitter_AQFP splitterN45ton332n333_( clk_4 , buf_splitterN45ton216n333_splitterN45ton332n333_1 , 0 , splitterN45ton332n333 );
splitter_AQFP splitterN49ton141n338_( clk_3 , N49 , 0 , splitterN49ton141n338 );
splitter_AQFP splitterN49ton42n338_( clk_5 , splitterN49ton141n338 , 0 , splitterN49ton42n338 );
splitter_AQFP splitterN49ton337n338_( clk_4 , buf_splitterN49ton42n338_splitterN49ton337n338_1 , 0 , splitterN49ton337n338 );
splitter_AQFP splitterN5ton186n288_( clk_2 , N5 , 0 , splitterN5ton186n288 );
splitter_AQFP splitterN5ton187n288_( clk_3 , splitterN5ton186n288 , 0 , splitterN5ton187n288 );
splitter_AQFP splitterN5ton287n288_( clk_4 , buf_splitterN5ton187n288_splitterN5ton287n288_1 , 0 , splitterN5ton287n288 );
splitter_AQFP splitterN53ton141n342_( clk_3 , N53 , 0 , splitterN53ton141n342 );
splitter_AQFP splitterN53ton182n342_( clk_5 , splitterN53ton141n342 , 0 , splitterN53ton182n342 );
splitter_AQFP splitterN53ton341n342_( clk_4 , buf_splitterN53ton182n342_splitterN53ton341n342_1 , 0 , splitterN53ton341n342 );
splitter_AQFP splitterN57ton138n346_( clk_3 , N57 , 0 , splitterN57ton138n346 );
splitter_AQFP splitterN57ton155n346_( clk_5 , splitterN57ton138n346 , 0 , splitterN57ton155n346 );
splitter_AQFP splitterN57ton345n346_( clk_4 , buf_splitterN57ton155n346_splitterN57ton345n346_1 , 0 , splitterN57ton345n346 );
splitter_AQFP splitterN61ton138n350_( clk_3 , N61 , 0 , splitterN61ton138n350 );
splitter_AQFP splitterN61ton216n350_( clk_5 , splitterN61ton138n350 , 0 , splitterN61ton216n350 );
splitter_AQFP splitterN61ton349n350_( clk_4 , buf_splitterN61ton216n350_splitterN61ton349n350_1 , 0 , splitterN61ton349n350 );
splitter_AQFP splitterN65ton245n363_( clk_2 , N65 , 0 , splitterN65ton245n363 );
splitter_AQFP splitterN65ton59n363_( clk_3 , splitterN65ton245n363 , 0 , splitterN65ton59n363 );
splitter_AQFP splitterN65ton362n363_( clk_2 , buf_splitterN65ton59n363_splitterN65ton362n363_1 , 0 , splitterN65ton362n363 );
splitter_AQFP splitterN69ton264n367_( clk_2 , N69 , 0 , splitterN69ton264n367 );
splitter_AQFP splitterN69ton59n367_( clk_3 , splitterN69ton264n367 , 0 , splitterN69ton59n367 );
splitter_AQFP splitterN69ton366n367_( clk_2 , buf_splitterN69ton59n367_splitterN69ton366n367_1 , 0 , splitterN69ton366n367 );
splitter_AQFP splitterN73ton55n371_( clk_2 , N73 , 0 , splitterN73ton55n371 );
splitter_AQFP splitterN73ton56n371_( clk_3 , splitterN73ton55n371 , 0 , splitterN73ton56n371 );
splitter_AQFP splitterN73ton370n371_( clk_2 , buf_splitterN73ton56n371_splitterN73ton370n371_1 , 0 , splitterN73ton370n371 );
splitter_AQFP splitterN77ton120n375_( clk_2 , N77 , 0 , splitterN77ton120n375 );
splitter_AQFP splitterN77ton56n375_( clk_3 , splitterN77ton120n375 , 0 , splitterN77ton56n375 );
splitter_AQFP splitterN77ton374n375_( clk_2 , buf_splitterN77ton56n375_splitterN77ton374n375_1 , 0 , splitterN77ton374n375 );
splitter_AQFP splitterN81ton245n381_( clk_2 , N81 , 0 , splitterN81ton245n381 );
splitter_AQFP splitterN81ton68n381_( clk_3 , splitterN81ton245n381 , 0 , splitterN81ton68n381 );
splitter_AQFP splitterN81ton380n381_( clk_2 , buf_splitterN81ton68n381_splitterN81ton380n381_1 , 0 , splitterN81ton380n381 );
splitter_AQFP splitterN85ton264n385_( clk_2 , N85 , 0 , splitterN85ton264n385 );
splitter_AQFP splitterN85ton68n385_( clk_3 , splitterN85ton264n385 , 0 , splitterN85ton68n385 );
splitter_AQFP splitterN85ton384n385_( clk_2 , buf_splitterN85ton68n385_splitterN85ton384n385_1 , 0 , splitterN85ton384n385 );
splitter_AQFP splitterN89ton64n389_( clk_2 , N89 , 0 , splitterN89ton64n389 );
splitter_AQFP splitterN89ton65n389_( clk_3 , splitterN89ton64n389 , 0 , splitterN89ton65n389 );
splitter_AQFP splitterN89ton388n389_( clk_2 , buf_splitterN89ton65n389_splitterN89ton388n389_1 , 0 , splitterN89ton388n389 );
splitter_AQFP splitterN9ton92n292_( clk_3 , N9 , 0 , splitterN9ton92n292 );
splitter_AQFP splitterN9ton158n292_( clk_5 , splitterN9ton92n292 , 0 , splitterN9ton158n292 );
splitter_AQFP splitterN9ton291n292_( clk_4 , buf_splitterN9ton158n292_splitterN9ton291n292_1 , 0 , splitterN9ton291n292 );
splitter_AQFP splitterN93ton120n393_( clk_2 , N93 , 0 , splitterN93ton120n393 );
splitter_AQFP splitterN93ton65n393_( clk_3 , splitterN93ton120n393 , 0 , splitterN93ton65n393 );
splitter_AQFP splitterN93ton392n393_( clk_2 , buf_splitterN93ton65n393_splitterN93ton392n393_1 , 0 , splitterN93ton392n393 );
splitter_AQFP splitterN97ton170n398_( clk_3 , N97 , 0 , splitterN97ton170n398 );
splitter_AQFP splitterN97ton241n398_( clk_5 , splitterN97ton170n398 , 0 , splitterN97ton241n398 );
splitter_AQFP splitterN97ton397n398_( clk_2 , buf_splitterN97ton241n398_splitterN97ton397n398_1 , 0 , splitterN97ton397n398 );
splitter_AQFP splitterfromn44_( clk_8 , n44 , 0 , splitterfromn44 );
splitter_AQFP splitterfromn45_( clk_5 , n45 , 0 , splitterfromn45 );
splitter_AQFP splitterfromn48_( clk_6 , n48 , 0 , splitterfromn48 );
splitter_AQFP splitterfromn51_( clk_1 , n51 , 0 , splitterfromn51 );
splitter_AQFP splitterfromn54_( clk_4 , n54 , 0 , splitterfromn54 );
splitter_AQFP splitterfromn57_( clk_6 , n57 , 0 , splitterfromn57 );
splitter_AQFP splitterfromn60_( clk_6 , n60 , 0 , splitterfromn60 );
splitter_AQFP splittern63ton176n74_( clk_1 , n63 , 0 , splittern63ton176n74 );
splitter_AQFP splitterfromn66_( clk_6 , n66 , 0 , splitterfromn66 );
splitter_AQFP splitterfromn69_( clk_6 , n69 , 0 , splitterfromn69 );
splitter_AQFP splittern72ton73n229_( clk_1 , n72 , 0 , splittern72ton73n229 );
splitter_AQFP splitterfromn75_( clk_4 , n75 , 0 , splitterfromn75 );
splitter_AQFP splittern78ton210n336_( clk_7 , n78 , 0 , splittern78ton210n336 );
splitter_AQFP splittern78ton238n336_( clk_1 , splittern78ton210n336 , 0 , splittern78ton238n336 );
splitter_AQFP splittern78ton282n336_( clk_2 , buf_splittern78ton238n336_splittern78ton282n336_1 , 0 , splittern78ton282n336 );
splitter_AQFP splitterfromn79_( clk_8 , n79 , 0 , splitterfromn79 );
splitter_AQFP splitterfromn82_( clk_6 , n82 , 0 , splitterfromn82 );
splitter_AQFP splitterfromn85_( clk_6 , n85 , 0 , splitterfromn85 );
splitter_AQFP splitterfromn88_( clk_1 , n88 , 0 , splitterfromn88 );
splitter_AQFP splitterfromn91_( clk_4 , n91 , 0 , splitterfromn91 );
splitter_AQFP splitterfromn94_( clk_6 , n94 , 0 , splitterfromn94 );
splitter_AQFP splitterfromn97_( clk_6 , n97 , 0 , splitterfromn97 );
splitter_AQFP splittern100ton110n255_( clk_1 , n100 , 0 , splittern100ton110n255 );
splitter_AQFP splitterfromn103_( clk_6 , n103 , 0 , splitterfromn103 );
splitter_AQFP splitterfromn106_( clk_6 , n106 , 0 , splitterfromn106 );
splitter_AQFP splittern109ton110n274_( clk_1 , n109 , 0 , splittern109ton110n274 );
splitter_AQFP splitterfromn112_( clk_4 , n112 , 0 , splitterfromn112 );
splitter_AQFP splittern115ton153n421_( clk_7 , n115 , 0 , splittern115ton153n421 );
splitter_AQFP splittern115ton353n421_( clk_1 , splittern115ton153n421 , 0 , splittern115ton353n421 );
splitter_AQFP splittern115ton369n421_( clk_8 , buf_splittern115ton353n421_splittern115ton369n421_1 , 0 , splittern115ton369n421 );
splitter_AQFP splitterfromn116_( clk_7 , buf_n116_splitterfromn116_1 , 0 , splitterfromn116 );
splitter_AQFP splitterfromn119_( clk_5 , n119 , 0 , splitterfromn119 );
splitter_AQFP splitterfromn122_( clk_5 , n122 , 0 , splitterfromn122 );
splitter_AQFP splitterfromn125_( clk_8 , n125 , 0 , splitterfromn125 );
splitter_AQFP splitterfromn128_( clk_4 , n128 , 0 , splitterfromn128 );
splitter_AQFP splitterfromn131_( clk_6 , n131 , 0 , splitterfromn131 );
splitter_AQFP splitterfromn134_( clk_5 , n134 , 0 , splitterfromn134 );
splitter_AQFP splittern137ton147n255_( clk_1 , n137 , 0 , splittern137ton147n255 );
splitter_AQFP splitterfromn140_( clk_6 , n140 , 0 , splitterfromn140 );
splitter_AQFP splitterfromn143_( clk_6 , n143 , 0 , splitterfromn143 );
splitter_AQFP splittern146ton147n274_( clk_1 , n146 , 0 , splittern146ton147n274 );
splitter_AQFP splitterfromn149_( clk_4 , n149 , 0 , splitterfromn149 );
splitter_AQFP splittern152ton153n425_( clk_7 , n152 , 0 , splittern152ton153n425 );
splitter_AQFP splittern152ton353n425_( clk_1 , splittern152ton153n425 , 0 , splittern152ton353n425 );
splitter_AQFP splittern152ton373n425_( clk_8 , buf_splittern152ton353n425_splittern152ton373n425_1 , 0 , splittern152ton373n425 );
splitter_AQFP splittern153ton355n318_( clk_1 , n153 , 0 , splittern153ton355n318 );
splitter_AQFP splittern153ton281n318_( clk_8 , buf_splittern153ton355n318_splittern153ton281n318_1 , 0 , splittern153ton281n318 );
splitter_AQFP splitterfromn154_( clk_2 , buf_n154_splitterfromn154_1 , 0 , splitterfromn154 );
splitter_AQFP splitterfromn157_( clk_8 , n157 , 0 , splitterfromn157 );
splitter_AQFP splitterfromn160_( clk_8 , n160 , 0 , splitterfromn160 );
splitter_AQFP splitterfromn163_( clk_3 , n163 , 0 , splitterfromn163 );
splitter_AQFP splitterfromn166_( clk_6 , n166 , 0 , splitterfromn166 );
splitter_AQFP splitterfromn169_( clk_6 , n169 , 0 , splitterfromn169 );
splitter_AQFP splitterfromn172_( clk_6 , n172 , 0 , splitterfromn172 );
splitter_AQFP splittern175ton176n205_( clk_1 , n175 , 0 , splittern175ton176n205 );
splitter_AQFP splitterfromn178_( clk_6 , n178 , 0 , splitterfromn178 );
splitter_AQFP splittern181ton211n344_( clk_1 , n181 , 0 , splittern181ton211n344 );
splitter_AQFP splittern181ton236n344_( clk_2 , splittern181ton211n344 , 0 , splittern181ton236n344 );
splitter_AQFP splittern181ton290n344_( clk_2 , buf_splittern181ton236n344_splittern181ton290n344_1 , 0 , splittern181ton290n344 );
splitter_AQFP splitterfromn184_( clk_1 , n184 , 0 , splitterfromn184 );
splitter_AQFP splitterfromn185_( clk_5 , n185 , 0 , splitterfromn185 );
splitter_AQFP splitterfromn188_( clk_6 , n188 , 0 , splitterfromn188 );
splitter_AQFP splitterfromn191_( clk_1 , n191 , 0 , splitterfromn191 );
splitter_AQFP splitterfromn194_( clk_4 , n194 , 0 , splitterfromn194 );
splitter_AQFP splitterfromn197_( clk_6 , n197 , 0 , splitterfromn197 );
splitter_AQFP splitterfromn200_( clk_6 , n200 , 0 , splitterfromn200 );
splitter_AQFP splittern203ton204n229_( clk_1 , n203 , 0 , splittern203ton204n229 );
splitter_AQFP splitterfromn206_( clk_4 , n206 , 0 , splitterfromn206 );
splitter_AQFP splittern209ton210n340_( clk_7 , n209 , 0 , splittern209ton210n340 );
splitter_AQFP splittern209ton238n340_( clk_2 , buf_splittern209ton210n340_splittern209ton238n340_1 , 0 , splittern209ton238n340 );
splitter_AQFP splittern209ton286n340_( clk_2 , buf_splittern209ton238n340_splittern209ton286n340_1 , 0 , splittern209ton286n340 );
splitter_AQFP splitterfromn210_( clk_1 , n210 , 0 , splitterfromn210 );
splitter_AQFP splitterfromn211_( clk_3 , n211 , 0 , splitterfromn211 );
splitter_AQFP splitterfromn212_( clk_1 , n212 , 0 , splitterfromn212 );
splitter_AQFP splitterfromn213_( clk_3 , n213 , 0 , splitterfromn213 );
splitter_AQFP splitterfromn215_( clk_2 , buf_n215_splitterfromn215_1 , 0 , splitterfromn215 );
splitter_AQFP splitterfromn218_( clk_8 , n218 , 0 , splitterfromn218 );
splitter_AQFP splitterfromn221_( clk_8 , n221 , 0 , splitterfromn221 );
splitter_AQFP splitterfromn224_( clk_3 , n224 , 0 , splitterfromn224 );
splitter_AQFP splitterfromn227_( clk_6 , n227 , 0 , splitterfromn227 );
splitter_AQFP splitterfromn230_( clk_6 , n230 , 0 , splitterfromn230 );
splitter_AQFP splittern233ton235n348_( clk_1 , n233 , 0 , splittern233ton235n348 );
splitter_AQFP splittern233ton236n348_( clk_2 , splittern233ton235n348 , 0 , splittern233ton236n348 );
splitter_AQFP splittern233ton234n348_( clk_4 , splittern233ton236n348 , 0 , splittern233ton234n348 );
splitter_AQFP splittern233ton294n348_( clk_2 , buf_splittern233ton234n348_splittern233ton294n348_1 , 0 , splittern233ton294n348 );
splitter_AQFP splitterfromn235_( clk_3 , n235 , 0 , splitterfromn235 );
splitter_AQFP splitterfromn240_( clk_7 , n240 , 0 , splitterfromn240 );
splitter_AQFP splitterfromn243_( clk_8 , n243 , 0 , splitterfromn243 );
splitter_AQFP splitterfromn244_( clk_5 , n244 , 0 , splitterfromn244 );
splitter_AQFP splitterfromn247_( clk_5 , n247 , 0 , splitterfromn247 );
splitter_AQFP splitterfromn250_( clk_8 , n250 , 0 , splitterfromn250 );
splitter_AQFP splitterfromn253_( clk_3 , n253 , 0 , splitterfromn253 );
splitter_AQFP splitterfromn256_( clk_4 , n256 , 0 , splitterfromn256 );
splitter_AQFP splittern259ton279n413_( clk_7 , n259 , 0 , splittern259ton279n413 );
splitter_AQFP splittern259ton356n413_( clk_1 , splittern259ton279n413 , 0 , splittern259ton356n413 );
splitter_AQFP splittern259ton361n413_( clk_8 , buf_splittern259ton356n413_splittern259ton361n413_1 , 0 , splittern259ton361n413 );
splitter_AQFP splitterfromn262_( clk_8 , n262 , 0 , splitterfromn262 );
splitter_AQFP splitterfromn263_( clk_4 , n263 , 0 , splitterfromn263 );
splitter_AQFP splitterfromn266_( clk_5 , n266 , 0 , splitterfromn266 );
splitter_AQFP splitterfromn269_( clk_8 , n269 , 0 , splitterfromn269 );
splitter_AQFP splitterfromn272_( clk_4 , n272 , 0 , splitterfromn272 );
splitter_AQFP splitterfromn275_( clk_4 , n275 , 0 , splitterfromn275 );
splitter_AQFP splittern278ton279n417_( clk_7 , n278 , 0 , splittern278ton279n417 );
splitter_AQFP splittern278ton356n417_( clk_1 , splittern278ton279n417 , 0 , splittern278ton356n417 );
splitter_AQFP splittern278ton365n417_( clk_8 , buf_splittern278ton356n417_splittern278ton365n417_1 , 0 , splittern278ton365n417 );
splitter_AQFP splitterfromn279_( clk_1 , n279 , 0 , splitterfromn279 );
splitter_AQFP splitterfromn280_( clk_1 , n280 , 0 , splitterfromn280 );
splitter_AQFP splittern281ton282n294_( clk_3 , n281 , 0 , splittern281ton282n294 );
splitter_AQFP splitterfromn282_( clk_5 , n282 , 0 , splitterfromn282 );
splitter_AQFP splitterfromn286_( clk_5 , n286 , 0 , splitterfromn286 );
splitter_AQFP splitterfromn290_( clk_5 , n290 , 0 , splitterfromn290 );
splitter_AQFP splitterfromn294_( clk_5 , n294 , 0 , splitterfromn294 );
splitter_AQFP splittern298ton355n335_( clk_1 , n298 , 0 , splittern298ton355n335 );
splitter_AQFP splittern298ton299n335_( clk_8 , buf_splittern298ton355n335_splittern298ton299n335_1 , 0 , splittern298ton299n335 );
splitter_AQFP splittern299ton300n312_( clk_3 , n299 , 0 , splittern299ton300n312 );
splitter_AQFP splitterfromn300_( clk_5 , n300 , 0 , splitterfromn300 );
splitter_AQFP splitterfromn304_( clk_5 , n304 , 0 , splitterfromn304 );
splitter_AQFP splitterfromn308_( clk_5 , n308 , 0 , splitterfromn308 );
splitter_AQFP splitterfromn312_( clk_5 , n312 , 0 , splitterfromn312 );
splitter_AQFP splitterfromn316_( clk_1 , n316 , 0 , splitterfromn316 );
splitter_AQFP splitterfromn317_( clk_1 , n317 , 0 , splitterfromn317 );
splitter_AQFP splittern318ton319n331_( clk_3 , n318 , 0 , splittern318ton319n331 );
splitter_AQFP splitterfromn319_( clk_5 , n319 , 0 , splitterfromn319 );
splitter_AQFP splitterfromn323_( clk_5 , n323 , 0 , splitterfromn323 );
splitter_AQFP splitterfromn327_( clk_5 , n327 , 0 , splitterfromn327 );
splitter_AQFP splitterfromn331_( clk_5 , n331 , 0 , splitterfromn331 );
splitter_AQFP splittern335ton336n348_( clk_3 , n335 , 0 , splittern335ton336n348 );
splitter_AQFP splitterfromn336_( clk_5 , n336 , 0 , splitterfromn336 );
splitter_AQFP splitterfromn340_( clk_5 , n340 , 0 , splitterfromn340 );
splitter_AQFP splitterfromn344_( clk_5 , n344 , 0 , splitterfromn344 );
splitter_AQFP splitterfromn348_( clk_5 , n348 , 0 , splitterfromn348 );
splitter_AQFP splitterfromn358_( clk_5 , n358 , 0 , splitterfromn358 );
splitter_AQFP splitterfromn359_( clk_7 , n359 , 0 , splitterfromn359 );
splitter_AQFP splittern360ton361n373_( clk_1 , n360 , 0 , splittern360ton361n373 );
splitter_AQFP splitterfromn361_( clk_3 , n361 , 0 , splitterfromn361 );
splitter_AQFP splitterfromn365_( clk_3 , n365 , 0 , splitterfromn365 );
splitter_AQFP splitterfromn369_( clk_3 , n369 , 0 , splitterfromn369 );
splitter_AQFP splitterfromn373_( clk_3 , n373 , 0 , splitterfromn373 );
splitter_AQFP splitterfromn377_( clk_7 , n377 , 0 , splitterfromn377 );
splitter_AQFP splittern378ton379n391_( clk_1 , n378 , 0 , splittern378ton379n391 );
splitter_AQFP splitterfromn379_( clk_3 , n379 , 0 , splitterfromn379 );
splitter_AQFP splitterfromn383_( clk_3 , n383 , 0 , splitterfromn383 );
splitter_AQFP splitterfromn387_( clk_3 , n387 , 0 , splitterfromn387 );
splitter_AQFP splitterfromn391_( clk_3 , n391 , 0 , splitterfromn391 );
splitter_AQFP splittern395ton396n408_( clk_1 , n395 , 0 , splittern395ton396n408 );
splitter_AQFP splitterfromn396_( clk_3 , n396 , 0 , splitterfromn396 );
splitter_AQFP splitterfromn400_( clk_3 , n400 , 0 , splitterfromn400 );
splitter_AQFP splitterfromn404_( clk_3 , n404 , 0 , splitterfromn404 );
splitter_AQFP splitterfromn408_( clk_3 , n408 , 0 , splitterfromn408 );
splitter_AQFP splittern412ton413n425_( clk_1 , n412 , 0 , splittern412ton413n425 );
splitter_AQFP splitterfromn413_( clk_3 , n413 , 0 , splitterfromn413 );
splitter_AQFP splitterfromn417_( clk_3 , n417 , 0 , splitterfromn417 );
splitter_AQFP splitterfromn421_( clk_3 , n421 , 0 , splitterfromn421 );
splitter_AQFP splitterfromn425_( clk_3 , n425 , 0 , splitterfromn425 );

endmodule