module top( clk_1 , clk_2 , clk_3 , clk_4 , clk_5 , clk_6 , clk_7 , clk_8 , G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G4 , G5 , G6 , G7 , G8 , G9 , G1884 , G1885 , G1886 , G1887 , G1888 , G1889 , G1890 , G1891 , G1892 , G1893 , G1894 , G1895 , G1896 , G1897 , G1898 , G1899 , G1900 , G1901 , G1902 , G1903 , G1904 , G1905 , G1906 , G1907 , G1908 );

input G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G4 , G5 , G6 , G7 , G8 , G9 ;
output G1884 , G1885 , G1886 , G1887 , G1888 , G1889 , G1890 , G1891 , G1892 , G1893 , G1894 , G1895 , G1896 , G1897 , G1898 , G1899 , G1900 , G1901 , G1902 , G1903 , G1904 , G1905 , G1906 , G1907 , G1908 ;
wire n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , buf_G1_splitterG1ton207n91_1 , buf_G1_splitterG1ton207n91_2 , buf_G12_splitterG12ton163n83_1 , buf_G16_splitterG16ton106n65_1 , buf_G16_splitterG16ton106n65_2 , buf_G17_splitterfromG17_1 , buf_G18_splitterfromG18_1 , buf_G19_splitterfromG19_1 , buf_G19_splitterfromG19_2 , buf_G20_splitterfromG20_1 , buf_G22_splitterfromG22_1 , buf_G24_splitterG24ton200n88_1 , buf_G25_splitterG25ton193n281_1 , buf_G25_splitterG25ton193n281_2 , buf_G25_splitterG25ton193n281_3 , buf_G25_splitterG25ton193n281_4 , buf_G25_splitterG25ton193n281_5 , buf_G25_splitterG25ton193n281_6 , buf_G25_splitterG25ton193n281_7 , buf_G25_splitterG25ton193n281_8 , buf_G25_splitterG25ton193n281_9 , buf_G26_splitterG26ton100n320_1 , buf_G26_splitterG26ton100n320_2 , buf_G26_splitterG26ton100n320_3 , buf_G26_splitterG26ton100n320_4 , buf_G26_splitterG26ton100n320_5 , buf_G26_splitterG26ton100n320_6 , buf_G26_splitterG26ton100n320_7 , buf_G27_splitterG27ton153n287_1 , buf_G27_splitterG27ton153n287_2 , buf_G27_splitterG27ton153n287_3 , buf_G27_splitterG27ton153n287_4 , buf_G27_splitterG27ton153n287_5 , buf_G27_splitterG27ton153n287_6 , buf_G27_splitterG27ton153n287_7 , buf_G28_splitterG28ton173n291_1 , buf_G28_splitterG28ton173n291_2 , buf_G28_splitterG28ton173n291_3 , buf_G28_splitterG28ton173n291_4 , buf_G28_splitterG28ton173n291_5 , buf_G28_splitterG28ton173n291_6 , buf_G28_splitterG28ton173n291_7 , buf_G28_splitterG28ton173n291_8 , buf_G29_splitterfromG29_1 , buf_G30_splitterfromG30_1 , buf_G32_splitterfromG32_1 , buf_G32_splitterfromG32_2 , buf_G32_splitterfromG32_3 , buf_n35_splittern35ton252n78_1 , buf_n35_splittern35ton252n78_2 , buf_n35_splittern35ton252n78_3 , buf_n57_splitterfromn57_1 , buf_n74_splittern74ton275n76_1 , buf_n122_splitterfromn122_1 , buf_n148_splitterfromn148_1 , buf_n148_splitterfromn148_2 , buf_n178_splittern178ton196n269_1 , buf_n178_splittern178ton196n269_2 , buf_n199_splitterfromn199_1 , buf_n199_splitterfromn199_2 , buf_n199_splitterfromn199_3 , buf_n200_splitterfromn200_1 , buf_n200_splitterfromn200_2 , buf_n202_n205_1 , buf_n203_splittern203ton204n321_1 , buf_n203_splittern203ton204n321_2 , buf_n203_splittern203ton204n321_3 , buf_n209_G1884_1 , buf_n209_G1884_2 , buf_n212_G1885_1 , buf_n214_n215_1 , buf_n215_G1886_1 , buf_n218_G1887_1 , buf_n218_G1887_2 , buf_n219_splitterfromn219_1 , buf_n219_splitterfromn219_2 , buf_n219_splitterfromn219_3 , buf_n219_splitterfromn219_4 , buf_n219_splitterfromn219_5 , buf_n221_splittern221ton222n254_1 , buf_n221_splittern221ton222n254_2 , buf_n225_G1888_1 , buf_n225_G1888_2 , buf_n225_G1888_3 , buf_n225_G1888_4 , buf_n226_n228_1 , buf_n228_G1889_1 , buf_n231_G1890_1 , buf_n231_G1890_2 , buf_n238_G1891_1 , buf_n238_G1891_2 , buf_n241_G1892_1 , buf_n241_G1892_2 , buf_n243_n244_1 , buf_n244_G1893_1 , buf_n247_G1894_1 , buf_n247_G1894_2 , buf_n247_G1894_3 , buf_n251_G1895_1 , buf_n251_G1895_2 , buf_n251_G1895_3 , buf_n251_G1895_4 , buf_n251_G1895_5 , buf_n257_G1896_1 , buf_n257_G1896_2 , buf_n260_G1897_1 , buf_n260_G1897_2 , buf_n260_G1897_3 , buf_n260_G1897_4 , buf_n263_G1898_1 , buf_n266_G1899_1 , buf_n266_G1899_2 , buf_n266_G1899_3 , buf_n273_n274_1 , buf_n273_n274_2 , buf_n273_n274_3 , buf_n274_G1900_1 , buf_n287_n288_1 , buf_n287_n288_2 , buf_n287_n288_3 , buf_n287_n288_4 , buf_n287_n288_5 , buf_n287_n288_6 , buf_n287_n288_7 , buf_n291_n292_1 , buf_n291_n292_2 , buf_n291_n292_3 , buf_n291_n292_4 , buf_n291_n292_5 , buf_n291_n292_6 , buf_n295_n296_1 , buf_n295_n296_2 , buf_n295_n296_3 , buf_n295_n296_4 , buf_n295_n296_5 , buf_n300_splitterfromn300_1 , buf_n300_splitterfromn300_2 , buf_n300_splitterfromn300_3 , buf_n300_splitterfromn300_4 , buf_n300_splitterfromn300_5 , buf_n308_n311_1 , buf_n308_n311_2 , buf_n309_n310_1 , buf_n311_splitterfromn311_1 , buf_n311_splitterfromn311_2 , buf_n311_splitterfromn311_3 , buf_n312_splitterfromn312_1 , buf_n312_splitterfromn312_2 , buf_n312_splitterfromn312_3 , buf_n312_splitterfromn312_4 , buf_splitterG1ton207n91_n207_1 , buf_splitterG1ton207n91_n207_2 , buf_splitterG1ton207n91_n207_3 , buf_splitterG1ton207n91_n207_4 , buf_splitterG1ton207n91_n207_5 , buf_splitterG1ton207n91_n207_6 , buf_splitterG1ton207n91_n207_7 , buf_splitterG1ton207n91_n207_8 , buf_splitterG1ton207n91_n207_9 , buf_splitterG1ton207n91_n207_10 , buf_splitterG1ton207n91_n207_11 , buf_splitterG1ton207n91_n207_12 , buf_splitterG1ton207n91_n208_1 , buf_splitterG1ton207n91_n208_2 , buf_splitterG1ton207n91_n208_3 , buf_splitterG1ton207n91_n208_4 , buf_splitterG1ton207n91_n208_5 , buf_splitterG1ton207n91_n208_6 , buf_splitterG1ton207n91_n208_7 , buf_splitterG1ton207n91_n208_8 , buf_splitterG1ton207n91_n208_9 , buf_splitterG1ton207n91_n208_10 , buf_splitterG1ton207n91_n208_11 , buf_splitterG1ton207n91_n208_12 , buf_splitterG10ton120n62_n120_1 , buf_splitterG10ton120n62_n121_1 , buf_splitterG10ton120n62_n223_1 , buf_splitterG10ton120n62_n223_2 , buf_splitterG10ton120n62_n223_3 , buf_splitterG10ton120n62_n223_4 , buf_splitterG10ton120n62_n223_5 , buf_splitterG10ton120n62_n223_6 , buf_splitterG10ton120n62_n223_7 , buf_splitterG10ton120n62_n223_8 , buf_splitterG10ton120n62_n223_9 , buf_splitterG10ton120n62_n223_10 , buf_splitterG10ton120n62_n223_11 , buf_splitterG10ton120n62_n223_12 , buf_splitterG10ton120n62_n223_13 , buf_splitterG10ton224n62_n224_1 , buf_splitterG10ton224n62_n224_2 , buf_splitterG10ton224n62_n224_3 , buf_splitterG10ton224n62_n224_4 , buf_splitterG10ton224n62_n224_5 , buf_splitterG10ton224n62_n224_6 , buf_splitterG10ton224n62_n224_7 , buf_splitterG10ton224n62_n224_8 , buf_splitterG10ton224n62_n224_9 , buf_splitterG10ton224n62_n224_10 , buf_splitterG10ton224n62_n224_11 , buf_splitterG10ton224n62_n224_12 , buf_splitterG10ton224n62_n224_13 , buf_splitterG11ton134n80_n255_1 , buf_splitterG11ton134n80_n255_2 , buf_splitterG11ton134n80_n255_3 , buf_splitterG11ton134n80_n255_4 , buf_splitterG11ton134n80_n255_5 , buf_splitterG11ton134n80_n255_6 , buf_splitterG11ton134n80_n255_7 , buf_splitterG11ton134n80_n255_8 , buf_splitterG11ton134n80_n255_9 , buf_splitterG11ton134n80_n255_10 , buf_splitterG11ton134n80_n255_11 , buf_splitterG11ton134n80_n255_12 , buf_splitterG11ton134n80_n255_13 , buf_splitterG11ton256n80_n256_1 , buf_splitterG11ton256n80_n256_2 , buf_splitterG11ton256n80_n256_3 , buf_splitterG11ton256n80_n256_4 , buf_splitterG11ton256n80_n256_5 , buf_splitterG11ton256n80_n256_6 , buf_splitterG11ton256n80_n256_7 , buf_splitterG11ton256n80_n256_8 , buf_splitterG11ton256n80_n256_9 , buf_splitterG11ton256n80_n256_10 , buf_splitterG11ton256n80_n256_11 , buf_splitterG11ton256n80_n256_12 , buf_splitterG11ton256n80_n256_13 , buf_splitterG12ton163n83_n258_1 , buf_splitterG12ton163n83_n258_2 , buf_splitterG12ton163n83_n258_3 , buf_splitterG12ton163n83_n258_4 , buf_splitterG12ton163n83_n258_5 , buf_splitterG12ton163n83_n258_6 , buf_splitterG12ton163n83_n258_7 , buf_splitterG12ton163n83_n258_8 , buf_splitterG12ton163n83_n258_9 , buf_splitterG12ton163n83_n258_10 , buf_splitterG12ton163n83_n258_11 , buf_splitterG12ton163n83_n258_12 , buf_splitterG12ton163n83_n258_13 , buf_splitterG12ton259n83_n259_1 , buf_splitterG12ton259n83_n259_2 , buf_splitterG12ton259n83_n259_3 , buf_splitterG12ton259n83_n259_4 , buf_splitterG12ton259n83_n259_5 , buf_splitterG12ton259n83_n259_6 , buf_splitterG12ton259n83_n259_7 , buf_splitterG12ton259n83_n259_8 , buf_splitterG12ton259n83_n259_9 , buf_splitterG12ton259n83_n259_10 , buf_splitterG12ton259n83_n259_11 , buf_splitterG12ton259n83_n259_12 , buf_splitterG13ton111n80_n111_1 , buf_splitterG13ton111n80_n111_2 , buf_splitterG13ton111n80_n112_1 , buf_splitterG13ton111n80_n112_2 , buf_splitterG13ton111n80_n261_1 , buf_splitterG13ton111n80_n261_2 , buf_splitterG13ton111n80_n261_3 , buf_splitterG13ton111n80_n261_4 , buf_splitterG13ton111n80_n261_5 , buf_splitterG13ton111n80_n261_6 , buf_splitterG13ton111n80_n261_7 , buf_splitterG13ton111n80_n261_8 , buf_splitterG13ton111n80_n261_9 , buf_splitterG13ton111n80_n261_10 , buf_splitterG13ton111n80_n261_11 , buf_splitterG13ton111n80_n261_12 , buf_splitterG13ton111n80_n261_13 , buf_splitterG13ton111n80_n261_14 , buf_splitterG13ton111n80_n261_15 , buf_splitterG13ton262n80_n262_1 , buf_splitterG13ton262n80_n262_2 , buf_splitterG13ton262n80_n262_3 , buf_splitterG13ton262n80_n262_4 , buf_splitterG13ton262n80_n262_5 , buf_splitterG13ton262n80_n262_6 , buf_splitterG13ton262n80_n262_7 , buf_splitterG13ton262n80_n262_8 , buf_splitterG13ton262n80_n262_9 , buf_splitterG13ton262n80_n262_10 , buf_splitterG13ton262n80_n262_11 , buf_splitterG13ton262n80_n262_12 , buf_splitterG13ton262n80_n262_13 , buf_splitterG13ton262n80_n262_14 , buf_splitterG14ton103n265_n180_1 , buf_splitterG14ton181n265_n264_1 , buf_splitterG14ton181n265_n264_2 , buf_splitterG14ton181n265_n264_3 , buf_splitterG14ton181n265_n264_4 , buf_splitterG14ton181n265_n264_5 , buf_splitterG14ton181n265_n264_6 , buf_splitterG14ton181n265_n264_7 , buf_splitterG14ton181n265_n264_8 , buf_splitterG14ton181n265_n264_9 , buf_splitterG14ton181n265_n264_10 , buf_splitterG14ton181n265_n264_11 , buf_splitterG14ton181n265_n264_12 , buf_splitterG14ton181n265_n264_13 , buf_splitterG14ton181n265_n265_1 , buf_splitterG14ton181n265_n265_2 , buf_splitterG14ton181n265_n265_3 , buf_splitterG14ton181n265_n265_4 , buf_splitterG14ton181n265_n265_5 , buf_splitterG14ton181n265_n265_6 , buf_splitterG14ton181n265_n265_7 , buf_splitterG14ton181n265_n265_8 , buf_splitterG14ton181n265_n265_9 , buf_splitterG14ton181n265_n265_10 , buf_splitterG14ton181n265_n265_11 , buf_splitterG14ton181n265_n265_12 , buf_splitterG14ton181n265_n265_13 , buf_splitterG15ton134n62_n226_1 , buf_splitterG15ton134n62_n226_2 , buf_splitterG15ton134n62_n226_3 , buf_splitterG15ton134n62_n226_4 , buf_splitterG15ton134n62_n226_5 , buf_splitterG15ton134n62_n226_6 , buf_splitterG15ton134n62_n226_7 , buf_splitterG15ton134n62_n226_8 , buf_splitterG15ton134n62_n226_9 , buf_splitterG15ton134n62_n226_10 , buf_splitterG15ton134n62_n226_11 , buf_splitterG15ton134n62_n226_12 , buf_splitterG15ton134n62_n226_13 , buf_splitterG15ton134n62_n226_14 , buf_splitterG15ton227n62_n227_1 , buf_splitterG15ton227n62_n227_2 , buf_splitterG15ton227n62_n227_3 , buf_splitterG15ton227n62_n227_4 , buf_splitterG15ton227n62_n227_5 , buf_splitterG15ton227n62_n227_6 , buf_splitterG15ton227n62_n227_7 , buf_splitterG15ton227n62_n227_8 , buf_splitterG15ton227n62_n227_9 , buf_splitterG15ton227n62_n227_10 , buf_splitterG15ton227n62_n227_11 , buf_splitterG15ton227n62_n227_12 , buf_splitterG15ton227n62_n227_13 , buf_splitterG15ton227n62_n227_14 , buf_splitterG16ton106n65_n229_1 , buf_splitterG16ton106n65_n229_2 , buf_splitterG16ton106n65_n229_3 , buf_splitterG16ton106n65_n229_4 , buf_splitterG16ton106n65_n229_5 , buf_splitterG16ton106n65_n229_6 , buf_splitterG16ton106n65_n229_7 , buf_splitterG16ton106n65_n229_8 , buf_splitterG16ton106n65_n229_9 , buf_splitterG16ton106n65_n229_10 , buf_splitterG16ton106n65_n229_11 , buf_splitterG16ton106n65_n229_12 , buf_splitterG16ton106n65_n229_13 , buf_splitterG16ton230n65_n230_1 , buf_splitterG16ton230n65_n230_2 , buf_splitterG16ton230n65_n230_3 , buf_splitterG16ton230n65_n230_4 , buf_splitterG16ton230n65_n230_5 , buf_splitterG16ton230n65_n230_6 , buf_splitterG16ton230n65_n230_7 , buf_splitterG16ton230n65_n230_8 , buf_splitterG16ton230n65_n230_9 , buf_splitterG16ton230n65_n230_10 , buf_splitterG16ton230n65_n230_11 , buf_splitterG16ton230n65_n230_12 , buf_splitterfromG17_n74_1 , buf_splitterfromG17_n74_2 , buf_splitterfromG17_n74_3 , buf_splitterfromG17_n74_4 , buf_splitterfromG17_n74_5 , buf_splitterfromG18_n35_1 , buf_splitterfromG18_n35_2 , buf_splitterfromG18_n35_3 , buf_splitterfromG19_n128_1 , buf_splitterfromG19_n128_2 , buf_splitterfromG19_n128_3 , buf_splitterfromG19_n128_4 , buf_splitterfromG19_n128_5 , buf_splitterG2ton146n46_n146_1 , buf_splitterG2ton146n46_n147_1 , buf_splitterG2ton146n46_n210_1 , buf_splitterG2ton146n46_n210_2 , buf_splitterG2ton146n46_n210_3 , buf_splitterG2ton146n46_n210_4 , buf_splitterG2ton146n46_n210_5 , buf_splitterG2ton146n46_n210_6 , buf_splitterG2ton146n46_n210_7 , buf_splitterG2ton146n46_n210_8 , buf_splitterG2ton146n46_n210_9 , buf_splitterG2ton146n46_n210_10 , buf_splitterG2ton146n46_n210_11 , buf_splitterG2ton146n46_n210_12 , buf_splitterG2ton146n46_n210_13 , buf_splitterG2ton146n46_n210_14 , buf_splitterG2ton211n46_n211_1 , buf_splitterG2ton211n46_n211_2 , buf_splitterG2ton211n46_n211_3 , buf_splitterG2ton211n46_n211_4 , buf_splitterG2ton211n46_n211_5 , buf_splitterG2ton211n46_n211_6 , buf_splitterG2ton211n46_n211_7 , buf_splitterG2ton211n46_n211_8 , buf_splitterG2ton211n46_n211_9 , buf_splitterG2ton211n46_n211_10 , buf_splitterG2ton211n46_n211_11 , buf_splitterG2ton211n46_n211_12 , buf_splitterG2ton211n46_n211_13 , buf_splitterG2ton211n46_n211_14 , buf_splitterfromG20_n178_1 , buf_splitterfromG20_n178_2 , buf_splitterfromG20_n178_3 , buf_splitterfromG20_n178_4 , buf_splitterfromG20_n178_5 , buf_splitterfromG20_n178_6 , buf_splitterG23ton109n200_n127_1 , buf_splitterG23ton109n200_n127_2 , buf_splitterG23ton109n200_n127_3 , buf_splitterG23ton109n200_n127_4 , buf_splitterG23ton109n200_n200_1 , buf_splitterG24ton200n88_n200_1 , buf_splitterG24ton200n88_n34_1 , buf_splitterG24ton200n88_n34_2 , buf_splitterG24ton200n88_n34_3 , buf_splitterG24ton200n88_n34_4 , buf_splitterG24ton200n88_n34_5 , buf_splitterG25ton193n281_n281_1 , buf_splitterG25ton193n281_n281_2 , buf_splitterG25ton193n281_n281_3 , buf_splitterG25ton193n281_n281_4 , buf_splitterG25ton193n281_n281_5 , buf_splitterG25ton193n281_n281_6 , buf_splitterG25ton193n281_n281_7 , buf_splitterG25ton193n281_n281_8 , buf_splitterG25ton193n281_n281_9 , buf_splitterG26ton100n320_n320_1 , buf_splitterG26ton100n320_n320_2 , buf_splitterG26ton100n320_n320_3 , buf_splitterG26ton100n320_n320_4 , buf_splitterG26ton100n320_n320_5 , buf_splitterG26ton100n320_n320_6 , buf_splitterG26ton100n320_n320_7 , buf_splitterG26ton100n320_n320_8 , buf_splitterG27ton153n287_n287_1 , buf_splitterG28ton173n291_n291_1 , buf_splitterfromG29_n199_1 , buf_splitterG3ton156n46_n213_1 , buf_splitterG3ton156n46_n213_2 , buf_splitterG3ton156n46_n213_3 , buf_splitterG3ton156n46_n213_4 , buf_splitterG3ton156n46_n213_5 , buf_splitterG3ton156n46_n213_6 , buf_splitterG3ton156n46_n213_7 , buf_splitterG3ton156n46_n213_8 , buf_splitterG3ton156n46_n213_9 , buf_splitterG3ton156n46_n213_10 , buf_splitterG3ton156n46_n213_11 , buf_splitterG3ton156n46_n213_12 , buf_splitterG3ton156n46_n213_13 , buf_splitterG3ton156n46_n213_14 , buf_splitterG3ton156n46_n213_15 , buf_splitterG3ton214n46_n214_1 , buf_splitterG3ton214n46_n214_2 , buf_splitterG3ton214n46_n214_3 , buf_splitterG3ton214n46_n214_4 , buf_splitterG3ton214n46_n214_5 , buf_splitterG3ton214n46_n214_6 , buf_splitterG3ton214n46_n214_7 , buf_splitterG3ton214n46_n214_8 , buf_splitterG3ton214n46_n214_9 , buf_splitterG3ton214n46_n214_10 , buf_splitterG3ton214n46_n214_11 , buf_splitterG3ton214n46_n214_12 , buf_splitterG3ton214n46_n214_13 , buf_splitterfromG30_n312_1 , buf_splitterG31ton126n127_n126_1 , buf_splitterG31ton126n127_n126_2 , buf_splitterG31ton152n201_n152_1 , buf_splitterG31ton152n201_n152_2 , buf_splitterG31ton152n201_n172_1 , buf_splitterG31ton152n201_n192_1 , buf_splitterG31ton152n201_n192_2 , buf_splitterG31ton276n291_n276_1 , buf_splitterG31ton276n291_n276_2 , buf_splitterG31ton276n291_n276_3 , buf_splitterG31ton276n291_n276_4 , buf_splitterG31ton276n291_n276_5 , buf_splitterG31ton276n291_n276_6 , buf_splitterG31ton276n291_n276_7 , buf_splitterG31ton276n291_n276_8 , buf_splitterG31ton276n291_n282_1 , buf_splitterG31ton276n291_n282_2 , buf_splitterG31ton276n291_n282_3 , buf_splitterG31ton276n291_n282_4 , buf_splitterG31ton276n291_n282_5 , buf_splitterG31ton276n291_n282_6 , buf_splitterG31ton276n291_n282_7 , buf_splitterG31ton276n291_n282_8 , buf_splitterG31ton295n99_n295_1 , buf_splitterG31ton295n99_n295_2 , buf_splitterG31ton295n99_n295_3 , buf_splitterG31ton295n99_n295_4 , buf_splitterG31ton295n99_n295_5 , buf_splitterG31ton295n99_n73_1 , buf_splitterG31ton295n99_n73_2 , buf_splitterG31ton295n99_n73_3 , buf_splitterG31ton295n99_n73_4 , buf_splitterG31ton295n99_n73_5 , buf_splitterG31ton295n99_n99_1 , buf_splitterG31ton295n99_n99_2 , buf_splitterG31ton295n99_n99_3 , buf_splitterfromG32_n268_1 , buf_splitterfromG32_n268_2 , buf_splitterfromG32_n268_3 , buf_splitterfromG32_n268_4 , buf_splitterfromG32_n268_5 , buf_splitterfromG32_n268_6 , buf_splitterfromG32_n268_7 , buf_splitterfromG32_n268_8 , buf_splitterfromG32_n268_9 , buf_splitterfromG32_n268_10 , buf_splitterfromG32_n268_11 , buf_splitterfromG32_n268_12 , buf_splitterfromG32_n268_13 , buf_splitterfromG32_n268_14 , buf_splitterG33ton109n88_n179_1 , buf_splitterG33ton199n273_n203_1 , buf_splitterG33ton199n273_n273_1 , buf_splitterG33ton199n273_n273_2 , buf_splitterG33ton199n273_n273_3 , buf_splitterG33ton199n273_n273_4 , buf_splitterG33ton199n273_n273_5 , buf_splitterG33ton199n273_n273_6 , buf_splitterG33ton199n273_n273_7 , buf_splitterG33ton199n273_n273_8 , buf_splitterG33ton199n273_n273_9 , buf_splitterG33ton199n273_n273_10 , buf_splitterG33ton199n273_n273_11 , buf_splitterG33ton304n88_n304_1 , buf_splitterG33ton304n88_n304_2 , buf_splitterG33ton304n88_n304_3 , buf_splitterG33ton304n88_n304_4 , buf_splitterG33ton304n88_n304_5 , buf_splitterG33ton304n88_n304_6 , buf_splitterG33ton304n88_n304_7 , buf_splitterG33ton304n88_n304_8 , buf_splitterG33ton304n88_n304_9 , buf_splitterG33ton304n88_n304_10 , buf_splitterG33ton304n88_n304_11 , buf_splitterG33ton304n88_n304_12 , buf_splitterG33ton304n88_n304_13 , buf_splitterG33ton304n88_n304_14 , buf_splitterG33ton304n88_n316_1 , buf_splitterG33ton304n88_n316_2 , buf_splitterG33ton304n88_n316_3 , buf_splitterG33ton304n88_n316_4 , buf_splitterG33ton304n88_n316_5 , buf_splitterG33ton304n88_n316_6 , buf_splitterG33ton304n88_n316_7 , buf_splitterG33ton304n88_n316_8 , buf_splitterG33ton304n88_n316_9 , buf_splitterG33ton304n88_n316_10 , buf_splitterG33ton304n88_n316_11 , buf_splitterG33ton304n88_n316_12 , buf_splitterG33ton304n88_n316_13 , buf_splitterG33ton304n88_n316_14 , buf_splitterG33ton304n88_n316_15 , buf_splitterG33ton304n88_n316_16 , buf_splitterG4ton216n43_n216_1 , buf_splitterG4ton216n43_n216_2 , buf_splitterG4ton216n43_n216_3 , buf_splitterG4ton216n43_n216_4 , buf_splitterG4ton216n43_n216_5 , buf_splitterG4ton216n43_n216_6 , buf_splitterG4ton216n43_n216_7 , buf_splitterG4ton216n43_n216_8 , buf_splitterG4ton216n43_n216_9 , buf_splitterG4ton216n43_n216_10 , buf_splitterG4ton216n43_n216_11 , buf_splitterG4ton216n43_n216_12 , buf_splitterG4ton216n43_n216_13 , buf_splitterG4ton216n43_n217_1 , buf_splitterG4ton216n43_n217_2 , buf_splitterG4ton216n43_n217_3 , buf_splitterG4ton216n43_n217_4 , buf_splitterG4ton216n43_n217_5 , buf_splitterG4ton216n43_n217_6 , buf_splitterG4ton216n43_n217_7 , buf_splitterG4ton216n43_n217_8 , buf_splitterG4ton216n43_n217_9 , buf_splitterG4ton216n43_n217_10 , buf_splitterG4ton216n43_n217_11 , buf_splitterG4ton216n43_n217_12 , buf_splitterG5ton143n40_n236_1 , buf_splitterG5ton143n40_n236_2 , buf_splitterG5ton143n40_n236_3 , buf_splitterG5ton143n40_n236_4 , buf_splitterG5ton143n40_n236_5 , buf_splitterG5ton143n40_n236_6 , buf_splitterG5ton143n40_n236_7 , buf_splitterG5ton143n40_n236_8 , buf_splitterG5ton143n40_n236_9 , buf_splitterG5ton143n40_n236_10 , buf_splitterG5ton143n40_n236_11 , buf_splitterG5ton143n40_n236_12 , buf_splitterG5ton143n40_n236_13 , buf_splitterG5ton237n40_n237_1 , buf_splitterG5ton237n40_n237_2 , buf_splitterG5ton237n40_n237_3 , buf_splitterG5ton237n40_n237_4 , buf_splitterG5ton237n40_n237_5 , buf_splitterG5ton237n40_n237_6 , buf_splitterG5ton237n40_n237_7 , buf_splitterG5ton237n40_n237_8 , buf_splitterG5ton237n40_n237_9 , buf_splitterG5ton237n40_n237_10 , buf_splitterG5ton237n40_n237_11 , buf_splitterG6ton156n37_n239_1 , buf_splitterG6ton156n37_n239_2 , buf_splitterG6ton156n37_n239_3 , buf_splitterG6ton156n37_n239_4 , buf_splitterG6ton156n37_n239_5 , buf_splitterG6ton156n37_n239_6 , buf_splitterG6ton156n37_n239_7 , buf_splitterG6ton156n37_n239_8 , buf_splitterG6ton156n37_n239_9 , buf_splitterG6ton156n37_n239_10 , buf_splitterG6ton156n37_n239_11 , buf_splitterG6ton156n37_n239_12 , buf_splitterG6ton156n37_n239_13 , buf_splitterG6ton156n37_n239_14 , buf_splitterG6ton240n37_n240_1 , buf_splitterG6ton240n37_n240_2 , buf_splitterG6ton240n37_n240_3 , buf_splitterG6ton240n37_n240_4 , buf_splitterG6ton240n37_n240_5 , buf_splitterG6ton240n37_n240_6 , buf_splitterG6ton240n37_n240_7 , buf_splitterG6ton240n37_n240_8 , buf_splitterG6ton240n37_n240_9 , buf_splitterG6ton240n37_n240_10 , buf_splitterG6ton240n37_n240_11 , buf_splitterG6ton240n37_n240_12 , buf_splitterG6ton240n37_n240_13 , buf_splitterG7ton117n37_n242_1 , buf_splitterG7ton117n37_n242_2 , buf_splitterG7ton117n37_n242_3 , buf_splitterG7ton117n37_n242_4 , buf_splitterG7ton117n37_n242_5 , buf_splitterG7ton117n37_n242_6 , buf_splitterG7ton117n37_n242_7 , buf_splitterG7ton117n37_n242_8 , buf_splitterG7ton117n37_n242_9 , buf_splitterG7ton117n37_n242_10 , buf_splitterG7ton117n37_n242_11 , buf_splitterG7ton117n37_n242_12 , buf_splitterG7ton117n37_n242_13 , buf_splitterG7ton117n37_n242_14 , buf_splitterG7ton243n37_n243_1 , buf_splitterG7ton243n37_n243_2 , buf_splitterG7ton243n37_n243_3 , buf_splitterG7ton243n37_n243_4 , buf_splitterG7ton243n37_n243_5 , buf_splitterG7ton243n37_n243_6 , buf_splitterG7ton243n37_n243_7 , buf_splitterG7ton243n37_n243_8 , buf_splitterG7ton243n37_n243_9 , buf_splitterG7ton243n37_n243_10 , buf_splitterG7ton243n37_n243_11 , buf_splitterG7ton243n37_n243_12 , buf_splitterG7ton243n37_n243_13 , buf_splitterG7ton243n37_n243_14 , buf_splitterG7ton243n37_n243_15 , buf_splitterG8ton245n43_n245_1 , buf_splitterG8ton245n43_n245_2 , buf_splitterG8ton245n43_n245_3 , buf_splitterG8ton245n43_n245_4 , buf_splitterG8ton245n43_n245_5 , buf_splitterG8ton245n43_n245_6 , buf_splitterG8ton245n43_n245_7 , buf_splitterG8ton245n43_n245_8 , buf_splitterG8ton245n43_n245_9 , buf_splitterG8ton245n43_n245_10 , buf_splitterG8ton245n43_n245_11 , buf_splitterG8ton245n43_n245_12 , buf_splitterG8ton245n43_n246_1 , buf_splitterG8ton245n43_n246_2 , buf_splitterG8ton245n43_n246_3 , buf_splitterG8ton245n43_n246_4 , buf_splitterG8ton245n43_n246_5 , buf_splitterG8ton245n43_n246_6 , buf_splitterG8ton245n43_n246_7 , buf_splitterG8ton245n43_n246_8 , buf_splitterG8ton245n43_n246_9 , buf_splitterG8ton245n43_n246_10 , buf_splitterG8ton245n43_n246_11 , buf_splitterG8ton245n43_n246_12 , buf_splitterG9ton103n59_n249_1 , buf_splitterG9ton103n59_n249_2 , buf_splitterG9ton103n59_n249_3 , buf_splitterG9ton103n59_n249_4 , buf_splitterG9ton103n59_n249_5 , buf_splitterG9ton103n59_n249_6 , buf_splitterG9ton103n59_n249_7 , buf_splitterG9ton103n59_n249_8 , buf_splitterG9ton103n59_n249_9 , buf_splitterG9ton103n59_n249_10 , buf_splitterG9ton103n59_n249_11 , buf_splitterG9ton103n59_n249_12 , buf_splitterG9ton103n59_n249_13 , buf_splitterG9ton250n59_n250_1 , buf_splitterG9ton250n59_n250_2 , buf_splitterG9ton250n59_n250_3 , buf_splitterG9ton250n59_n250_4 , buf_splitterG9ton250n59_n250_5 , buf_splitterG9ton250n59_n250_6 , buf_splitterG9ton250n59_n250_7 , buf_splitterG9ton250n59_n250_8 , buf_splitterG9ton250n59_n250_9 , buf_splitterG9ton250n59_n250_10 , buf_splitterG9ton250n59_n250_11 , buf_splitterfromn34_n74_1 , buf_splittern35ton252n78_n252_1 , buf_splittern35ton252n78_n252_2 , buf_splittern35ton252n78_n78_1 , buf_splittern41ton54n94_n54_1 , buf_splittern41ton54n94_n55_1 , buf_splittern50ton186n52_n186_1 , buf_splittern50ton186n52_n187_1 , buf_splittern66ton67n86_n67_1 , buf_splittern66ton67n86_n68_1 , buf_splitterfromn72_n277_1 , buf_splitterfromn72_n277_2 , buf_splitterfromn72_n277_3 , buf_splitterfromn72_n277_4 , buf_splitterfromn72_n277_5 , buf_splitterfromn72_n277_6 , buf_splitterfromn72_n277_7 , buf_splitterfromn72_n277_8 , buf_splitterfromn72_n277_9 , buf_splittern73ton278n76_n278_1 , buf_splittern73ton278n76_n278_2 , buf_splittern73ton278n76_n278_3 , buf_splittern73ton278n76_n278_4 , buf_splittern73ton278n76_n278_5 , buf_splittern73ton278n76_n278_6 , buf_splittern73ton278n76_n278_7 , buf_splittern74ton275n76_n275_1 , buf_splittern74ton275n76_n275_2 , buf_splittern74ton275n76_n275_3 , buf_splittern74ton275n76_n275_4 , buf_splittern74ton275n76_n275_5 , buf_splittern74ton275n76_n275_6 , buf_splittern74ton275n76_n275_7 , buf_splittern74ton275n76_n275_8 , buf_splittern77ton253n78_n253_1 , buf_splittern87ton189n97_n189_1 , buf_splittern87ton189n97_n190_1 , buf_splitterfromn98_n321_1 , buf_splitterfromn98_n321_2 , buf_splitterfromn98_n321_3 , buf_splitterfromn98_n321_4 , buf_splitterfromn98_n321_5 , buf_splitterfromn98_n321_6 , buf_splitterfromn98_n321_7 , buf_splitterfromn98_n321_8 , buf_splitterfromn98_n321_9 , buf_splitterfromn98_n321_10 , buf_splittern105ton106n309_n308_1 , buf_splittern105ton106n309_n308_2 , buf_splittern105ton106n309_n308_3 , buf_splittern105ton106n309_n309_1 , buf_splittern105ton106n309_n309_2 , buf_splittern105ton106n309_n309_3 , buf_splittern105ton106n309_n309_4 , buf_splitterfromn125_n297_1 , buf_splitterfromn125_n297_2 , buf_splitterfromn125_n297_3 , buf_splitterfromn125_n297_4 , buf_splitterfromn125_n297_5 , buf_splitterfromn125_n297_6 , buf_splitterfromn125_n297_7 , buf_splitterfromn125_n297_8 , buf_splitterfromn125_n297_9 , buf_splitterfromn125_n297_10 , buf_splittern128ton129n295_n295_1 , buf_splitterfromn151_n289_1 , buf_splitterfromn151_n289_2 , buf_splitterfromn151_n289_3 , buf_splitterfromn151_n289_4 , buf_splitterfromn151_n289_5 , buf_splitterfromn151_n289_6 , buf_splitterfromn151_n289_7 , buf_splitterfromn151_n289_8 , buf_splitterfromn151_n289_9 , buf_splitterfromn171_n293_1 , buf_splitterfromn171_n293_2 , buf_splitterfromn171_n293_3 , buf_splitterfromn171_n293_4 , buf_splitterfromn171_n293_5 , buf_splitterfromn171_n293_6 , buf_splitterfromn171_n293_7 , buf_splitterfromn171_n293_8 , buf_splitterfromn171_n293_9 , buf_splittern177ton197n272_n272_1 , buf_splitterfromn191_n283_1 , buf_splitterfromn191_n283_2 , buf_splitterfromn191_n283_3 , buf_splitterfromn191_n283_4 , buf_splitterfromn191_n283_5 , buf_splitterfromn191_n283_6 , buf_splitterfromn191_n283_7 , buf_splitterfromn191_n283_8 , buf_splitterfromn191_n283_9 , buf_splitterfromn191_n283_10 , buf_splittern192ton193n284_n284_1 , buf_splittern192ton193n284_n284_2 , buf_splittern192ton193n284_n284_3 , buf_splittern192ton193n284_n284_4 , buf_splittern192ton193n284_n284_5 , buf_splittern192ton193n284_n284_6 , buf_splittern192ton193n284_n284_7 , buf_splitterfromn200_n204_1 , buf_splittern203ton204n321_n279_1 , buf_splittern203ton204n321_n279_2 , buf_splittern203ton204n321_n279_3 , buf_splittern203ton204n321_n279_4 , buf_splittern203ton204n321_n279_5 , buf_splittern203ton204n321_n279_6 , buf_splittern203ton204n321_n279_7 , buf_splittern203ton204n321_n279_8 , buf_splittern203ton204n321_n279_9 , buf_splittern203ton204n321_n279_10 , buf_splittern203ton204n321_n279_11 , buf_splittern203ton204n321_n279_12 , buf_splittern203ton204n321_n279_13 , buf_splittern203ton204n321_n285_1 , buf_splittern203ton204n321_n285_2 , buf_splittern203ton204n321_n285_3 , buf_splittern203ton204n321_n285_4 , buf_splittern203ton204n321_n285_5 , buf_splittern203ton204n321_n285_6 , buf_splittern203ton204n321_n285_7 , buf_splittern203ton204n321_n285_8 , buf_splittern203ton204n321_n285_9 , buf_splittern203ton204n321_n285_10 , buf_splittern203ton204n321_n285_11 , buf_splittern203ton204n321_n285_12 , buf_splittern203ton204n321_n285_13 , buf_splittern203ton204n321_n285_14 , buf_splittern203ton290n321_n290_1 , buf_splittern203ton290n321_n294_1 , buf_splitterfromn205_n206_1 , buf_splitterfromn205_n206_2 , buf_splitterfromn205_n206_3 , buf_splitterfromn205_n206_4 , buf_splitterfromn205_n235_1 , buf_splitterfromn205_n235_2 , buf_splitterfromn205_n235_3 , buf_splitterfromn205_n235_4 , buf_splitterfromn205_n235_5 , buf_splitterfromn205_n235_6 , buf_splitterfromn219_n310_1 , buf_splittern221ton222n254_n222_1 , buf_splittern221ton222n254_n222_2 , buf_splittern221ton222n254_n248_1 , buf_splittern221ton222n254_n248_2 , buf_splittern221ton222n254_n254_1 , buf_splittern221ton222n254_n254_2 , buf_splitterfromn299_n305_1 , buf_splitterfromn299_n305_2 , buf_splitterfromn299_n305_3 , buf_splitterfromn299_n305_4 , buf_splitterfromn299_n305_5 , buf_splitterfromn299_n305_6 , buf_splitterfromn299_n305_7 , buf_splitterfromn299_n305_8 , buf_splitterfromn299_n306_1 , buf_splitterfromn299_n306_2 , buf_splitterfromn299_n306_3 , buf_splitterfromn299_n306_4 , buf_splitterfromn299_n306_5 , buf_splitterfromn299_n306_6 , buf_splitterfromn299_n306_7 , buf_splitterfromn299_n306_8 , buf_splitterfromn300_n301_1 , buf_splitterfromn300_n301_2 , buf_splitterfromn300_n301_3 , buf_splitterfromn300_n301_4 , buf_splitterfromn300_n301_5 , buf_splitterfromn300_n301_6 , buf_splitterfromn300_n301_7 , buf_splitterfromn300_n301_8 , buf_splitterfromn300_n301_9 , buf_splitterfromn300_n302_1 , buf_splitterfromn300_n302_2 , buf_splitterfromn300_n302_3 , buf_splitterfromn300_n302_4 , buf_splitterfromn300_n302_5 , buf_splitterfromn300_n302_6 , buf_splitterfromn300_n302_7 , buf_splitterfromn300_n302_8 , buf_splitterfromn300_n302_9 , buf_splitterfromn300_n302_10 , buf_splitterfromn311_n317_1 , buf_splitterfromn311_n317_2 , buf_splitterfromn311_n317_3 , buf_splitterfromn311_n318_1 , buf_splitterfromn311_n318_2 , buf_splitterfromn311_n318_3 , buf_splitterfromn311_n318_4 , buf_splitterfromn312_n313_1 , buf_splitterfromn312_n313_2 , buf_splitterfromn312_n313_3 , buf_splitterfromn312_n313_4 , buf_splitterfromn312_n313_5 , buf_splitterfromn312_n313_6 , buf_splitterfromn312_n313_7 , buf_splitterfromn312_n313_8 , buf_splitterfromn312_n313_9 , buf_splitterfromn312_n313_10 , buf_splitterfromn312_n314_1 , buf_splitterfromn312_n314_2 , buf_splitterfromn312_n314_3 , buf_splitterfromn312_n314_4 , buf_splitterfromn312_n314_5 , buf_splitterfromn312_n314_6 , buf_splitterfromn312_n314_7 , buf_splitterfromn312_n314_8 , buf_splitterfromn312_n314_9 , buf_splitterfromn312_n314_10 , buf_splitterfromn312_n314_11 , buf_splitterfromn312_n314_12 , splitterG1ton207n91 , splitterG1ton49n91 , splitterG10ton120n62 , splitterG10ton224n62 , splitterG11ton134n80 , splitterG11ton256n80 , splitterG12ton163n83 , splitterG12ton259n83 , splitterG13ton111n80 , splitterG13ton262n80 , splitterG14ton103n265 , splitterG14ton181n265 , splitterG15ton134n62 , splitterG15ton227n62 , splitterG16ton106n65 , splitterG16ton230n65 , splitterfromG17 , splitterfromG18 , splitterfromG19 , splitterG2ton146n46 , splitterG2ton211n46 , splitterfromG20 , splitterfromG21 , splitterfromG22 , splitterG23ton109n200 , splitterG24ton200n88 , splitterG25ton193n281 , splitterG26ton100n320 , splitterG27ton153n287 , splitterG28ton173n291 , splitterfromG29 , splitterG3ton156n46 , splitterG3ton214n46 , splitterfromG30 , splitterG31ton126n99 , splitterG31ton126n127 , splitterG31ton152n201 , splitterG31ton276n291 , splitterG31ton295n99 , splitterfromG32 , splitterG33ton109n88 , splitterG33ton199n273 , splitterG33ton304n88 , splitterG4ton117n43 , splitterG4ton180n181 , splitterG4ton216n43 , splitterG5ton143n40 , splitterG5ton237n40 , splitterG6ton156n37 , splitterG6ton240n37 , splitterG7ton117n37 , splitterG7ton243n37 , splitterG8ton143n43 , splitterG8ton159n160 , splitterG8ton245n43 , splitterG9ton103n59 , splitterG9ton250n59 , splitterfromn34 , splittern35ton252n78 , splitterfromn38 , splittern41ton54n94 , splitterfromn44 , splitterfromn47 , splittern50ton186n52 , splitterfromn53 , splittern56ton299n71 , splitterfromn57 , splitterfromn60 , splittern63ton163n65 , splittern66ton67n86 , splitterfromn69 , splitterfromn72 , splittern73ton278n76 , splittern74ton275n76 , splittern77ton253n78 , splitterfromn78 , splitterfromn81 , splitterfromn84 , splittern87ton189n97 , splittern87ton309n97 , splitterfromn88 , splitterfromn89 , splitterfromn92 , splitterfromn95 , splitterfromn98 , splitterfromn99 , splittern105ton106n309 , splittern108ton114n141 , splitterfromn109 , splitterfromn110 , splitterfromn113 , splitterfromn116 , splitterfromn119 , splitterfromn122 , splitterfromn125 , splitterfromn126 , splitterfromn127 , splittern128ton129n295 , splitterfromn133 , splitterfromn136 , splitterfromn139 , splitterfromn142 , splitterfromn145 , splitterfromn148 , splitterfromn151 , splitterfromn152 , splitterfromn158 , splitterfromn161 , splitterfromn162 , splitterfromn165 , splitterfromn168 , splitterfromn171 , splitterfromn172 , splittern177ton197n272 , splittern178ton196n269 , splitterfromn179 , splitterfromn182 , splitterfromn185 , splitterfromn188 , splitterfromn191 , splittern192ton193n284 , splittern195ton196n270 , splitterfromn197 , splitterfromn198 , splitterfromn199 , splitterfromn200 , splitterfromn201 , splittern203ton204n321 , splittern203ton290n321 , splitterfromn204 , splitterfromn205 , splittern206ton207n302 , splittern206ton208n210 , splittern206ton211n216 , splittern206ton217n302 , splitterfromn219 , splittern221ton222n254 , splittern222ton223n314 , splittern222ton226n229 , splittern222ton230n314 , splitterfromn234 , splittern235ton236n246 , splittern235ton239n240 , splittern235ton242n246 , splitterfromn248 , splittern254ton255n265 , splittern254ton258n259 , splittern254ton261n265 , splittern267ton268n320 , splittern267ton288n320 , splitterfromn275 , splitterfromn281 , splitterfromn299 , splitterfromn300 , splitterfromn304 , splitterfromn311 , splitterfromn312 , splitterfromn316 ;

PI_AQFP G1_( clk_1 , G1 );
PI_AQFP G10_( clk_1 , G10 );
PI_AQFP G11_( clk_1 , G11 );
PI_AQFP G12_( clk_1 , G12 );
PI_AQFP G13_( clk_1 , G13 );
PI_AQFP G14_( clk_1 , G14 );
PI_AQFP G15_( clk_1 , G15 );
PI_AQFP G16_( clk_1 , G16 );
PI_AQFP G17_( clk_1 , G17 );
PI_AQFP G18_( clk_1 , G18 );
PI_AQFP G19_( clk_1 , G19 );
PI_AQFP G2_( clk_1 , G2 );
PI_AQFP G20_( clk_1 , G20 );
PI_AQFP G21_( clk_1 , G21 );
PI_AQFP G22_( clk_1 , G22 );
PI_AQFP G23_( clk_1 , G23 );
PI_AQFP G24_( clk_1 , G24 );
PI_AQFP G25_( clk_1 , G25 );
PI_AQFP G26_( clk_1 , G26 );
PI_AQFP G27_( clk_1 , G27 );
PI_AQFP G28_( clk_1 , G28 );
PI_AQFP G29_( clk_1 , G29 );
PI_AQFP G3_( clk_1 , G3 );
PI_AQFP G30_( clk_1 , G30 );
PI_AQFP G31_( clk_1 , G31 );
PI_AQFP G32_( clk_1 , G32 );
PI_AQFP G33_( clk_1 , G33 );
PI_AQFP G4_( clk_1 , G4 );
PI_AQFP G5_( clk_1 , G5 );
PI_AQFP G6_( clk_1 , G6 );
PI_AQFP G7_( clk_1 , G7 );
PI_AQFP G8_( clk_1 , G8 );
PI_AQFP G9_( clk_1 , G9 );
or_AQFP n34_( clk_3 , buf_splitterG24ton200n88_n34_5 , splitterG31ton295n99 , 0 , 0 , n34 );
and_AQFP n35_( clk_5 , buf_splitterfromG18_n35_3 , splitterfromn34 , 0 , 0 , n35 );
or_AQFP n36_( clk_5 , splitterG6ton240n37 , splitterG7ton243n37 , 0 , 0 , n36 );
and_AQFP n37_( clk_5 , splitterG6ton240n37 , splitterG7ton243n37 , 0 , 0 , n37 );
and_AQFP n38_( clk_6 , n36 , n37 , 0 , 1 , n38 );
and_AQFP n39_( clk_8 , splitterG5ton237n40 , splitterfromn38 , 0 , 0 , n39 );
or_AQFP n40_( clk_8 , splitterG5ton237n40 , splitterfromn38 , 0 , 0 , n40 );
and_AQFP n41_( clk_1 , n39 , n40 , 1 , 0 , n41 );
or_AQFP n42_( clk_7 , splitterG4ton216n43 , splitterG8ton245n43 , 0 , 0 , n42 );
and_AQFP n43_( clk_7 , splitterG4ton216n43 , splitterG8ton245n43 , 0 , 0 , n43 );
and_AQFP n44_( clk_8 , n42 , n43 , 0 , 1 , n44 );
or_AQFP n45_( clk_4 , splitterG2ton211n46 , splitterG3ton214n46 , 0 , 0 , n45 );
and_AQFP n46_( clk_4 , splitterG2ton211n46 , splitterG3ton214n46 , 0 , 0 , n46 );
and_AQFP n47_( clk_5 , n45 , n46 , 0 , 1 , n47 );
and_AQFP n48_( clk_7 , splitterG1ton207n91 , splitterfromn47 , 0 , 0 , n48 );
or_AQFP n49_( clk_7 , splitterG1ton49n91 , splitterfromn47 , 0 , 0 , n49 );
and_AQFP n50_( clk_8 , n48 , n49 , 1 , 0 , n50 );
and_AQFP n51_( clk_2 , splitterfromn44 , splittern50ton186n52 , 1 , 0 , n51 );
and_AQFP n52_( clk_2 , splitterfromn44 , splittern50ton186n52 , 0 , 1 , n52 );
or_AQFP n53_( clk_3 , n51 , n52 , 0 , 0 , n53 );
or_AQFP n54_( clk_5 , buf_splittern41ton54n94_n54_1 , splitterfromn53 , 0 , 0 , n54 );
and_AQFP n55_( clk_5 , buf_splittern41ton54n94_n55_1 , splitterfromn53 , 0 , 0 , n55 );
and_AQFP n56_( clk_6 , n54 , n55 , 0 , 1 , n56 );
and_AQFP n57_( clk_5 , splitterfromG21 , splitterG33ton304n88 , 0 , 1 , n57 );
and_AQFP n58_( clk_1 , splitterG9ton250n59 , splitterfromn57 , 1 , 0 , n58 );
and_AQFP n59_( clk_1 , splitterG9ton250n59 , splitterfromn57 , 0 , 1 , n59 );
or_AQFP n60_( clk_2 , n58 , n59 , 0 , 0 , n60 );
and_AQFP n61_( clk_4 , splitterG10ton224n62 , splitterG15ton227n62 , 0 , 1 , n61 );
and_AQFP n62_( clk_4 , splitterG10ton224n62 , splitterG15ton227n62 , 1 , 0 , n62 );
or_AQFP n63_( clk_5 , n61 , n62 , 0 , 0 , n63 );
and_AQFP n64_( clk_7 , splitterG16ton230n65 , splittern63ton163n65 , 1 , 0 , n64 );
and_AQFP n65_( clk_7 , splitterG16ton230n65 , splittern63ton163n65 , 0 , 1 , n65 );
or_AQFP n66_( clk_8 , n64 , n65 , 0 , 0 , n66 );
and_AQFP n67_( clk_4 , splitterfromn60 , buf_splittern66ton67n86_n67_1 , 1 , 0 , n67 );
and_AQFP n68_( clk_4 , splitterfromn60 , buf_splittern66ton67n86_n68_1 , 0 , 1 , n68 );
or_AQFP n69_( clk_6 , n67 , n68 , 0 , 0 , n69 );
and_AQFP n70_( clk_8 , splittern56ton299n71 , splitterfromn69 , 0 , 1 , n70 );
and_AQFP n71_( clk_8 , splittern56ton299n71 , splitterfromn69 , 1 , 0 , n71 );
or_AQFP n72_( clk_1 , n70 , n71 , 0 , 0 , n72 );
or_AQFP n73_( clk_3 , buf_splitterG31ton295n99_n73_5 , splitterfromn72 , 0 , 0 , n73 );
and_AQFP n74_( clk_7 , buf_splitterfromG17_n74_5 , buf_splitterfromn34_n74_1 , 0 , 0 , n74 );
and_AQFP n75_( clk_5 , splittern73ton278n76 , splittern74ton275n76 , 0 , 1 , n75 );
and_AQFP n76_( clk_5 , splittern73ton278n76 , splittern74ton275n76 , 1 , 0 , n76 );
or_AQFP n77_( clk_6 , n75 , n76 , 0 , 0 , n77 );
and_AQFP n78_( clk_8 , buf_splittern35ton252n78_n78_1 , splittern77ton253n78 , 0 , 1 , n78 );
and_AQFP n79_( clk_4 , splitterG11ton256n80 , splitterG13ton262n80 , 1 , 0 , n79 );
and_AQFP n80_( clk_4 , splitterG11ton256n80 , splitterG13ton262n80 , 0 , 1 , n80 );
or_AQFP n81_( clk_5 , n79 , n80 , 0 , 0 , n81 );
and_AQFP n82_( clk_7 , splitterG12ton259n83 , splitterfromn81 , 0 , 1 , n82 );
and_AQFP n83_( clk_7 , splitterG12ton259n83 , splitterfromn81 , 1 , 0 , n83 );
or_AQFP n84_( clk_8 , n82 , n83 , 0 , 0 , n84 );
and_AQFP n85_( clk_2 , splittern66ton67n86 , splitterfromn84 , 1 , 0 , n85 );
and_AQFP n86_( clk_2 , splittern66ton67n86 , splitterfromn84 , 0 , 1 , n86 );
or_AQFP n87_( clk_3 , n85 , n86 , 0 , 0 , n87 );
or_AQFP n88_( clk_4 , splitterG24ton200n88 , splitterG33ton304n88 , 0 , 0 , n88 );
and_AQFP n89_( clk_6 , splitterfromG17 , splitterfromn88 , 0 , 1 , n89 );
and_AQFP n90_( clk_8 , splitterG1ton49n91 , splitterfromn89 , 1 , 0 , n90 );
and_AQFP n91_( clk_8 , splitterG1ton49n91 , splitterfromn89 , 0 , 1 , n91 );
or_AQFP n92_( clk_1 , n90 , n91 , 0 , 0 , n92 );
or_AQFP n93_( clk_3 , splittern41ton54n94 , splitterfromn92 , 0 , 0 , n93 );
and_AQFP n94_( clk_3 , splittern41ton54n94 , splitterfromn92 , 0 , 0 , n94 );
and_AQFP n95_( clk_4 , n93 , n94 , 0 , 1 , n95 );
or_AQFP n96_( clk_6 , splittern87ton309n97 , splitterfromn95 , 0 , 0 , n96 );
and_AQFP n97_( clk_6 , splittern87ton309n97 , splitterfromn95 , 0 , 0 , n97 );
and_AQFP n98_( clk_7 , n96 , n97 , 0 , 1 , n98 );
or_AQFP n99_( clk_1 , buf_splitterG31ton295n99_n99_3 , splitterfromn98 , 0 , 0 , n99 );
or_AQFP n100_( clk_3 , splitterG26ton100n320 , splitterfromn99 , 0 , 0 , n100 );
and_AQFP n101_( clk_3 , splitterG26ton100n320 , splitterfromn99 , 0 , 0 , n101 );
and_AQFP n102_( clk_4 , n100 , n101 , 0 , 1 , n102 );
and_AQFP n103_( clk_4 , splitterG14ton103n265 , splitterG9ton103n59 , 1 , 0 , n103 );
and_AQFP n104_( clk_4 , splitterG14ton103n265 , splitterG9ton103n59 , 0 , 1 , n104 );
or_AQFP n105_( clk_5 , n103 , n104 , 0 , 0 , n105 );
and_AQFP n106_( clk_7 , splitterG16ton106n65 , splittern105ton106n309 , 1 , 0 , n106 );
and_AQFP n107_( clk_7 , splitterG16ton106n65 , splittern105ton106n309 , 0 , 1 , n107 );
or_AQFP n108_( clk_1 , n106 , n107 , 0 , 0 , n108 );
or_AQFP n109_( clk_4 , splitterG23ton109n200 , splitterG33ton109n88 , 0 , 0 , n109 );
and_AQFP n110_( clk_6 , splitterfromG20 , splitterfromn109 , 0 , 1 , n110 );
and_AQFP n111_( clk_8 , buf_splitterG13ton111n80_n111_2 , splitterfromn110 , 1 , 0 , n111 );
and_AQFP n112_( clk_8 , buf_splitterG13ton111n80_n112_2 , splitterfromn110 , 0 , 1 , n112 );
or_AQFP n113_( clk_1 , n111 , n112 , 0 , 0 , n113 );
and_AQFP n114_( clk_3 , splittern108ton114n141 , splitterfromn113 , 1 , 0 , n114 );
and_AQFP n115_( clk_3 , splittern108ton114n141 , splitterfromn113 , 0 , 1 , n115 );
or_AQFP n116_( clk_4 , n114 , n115 , 0 , 0 , n116 );
and_AQFP n117_( clk_3 , splitterG4ton117n43 , splitterG7ton117n37 , 0 , 1 , n117 );
and_AQFP n118_( clk_3 , splitterG4ton117n43 , splitterG7ton117n37 , 1 , 0 , n118 );
or_AQFP n119_( clk_4 , n117 , n118 , 0 , 0 , n119 );
and_AQFP n120_( clk_6 , buf_splitterG10ton120n62_n120_1 , splitterfromn119 , 0 , 1 , n120 );
and_AQFP n121_( clk_6 , buf_splitterG10ton120n62_n121_1 , splitterfromn119 , 1 , 0 , n121 );
or_AQFP n122_( clk_8 , n120 , n121 , 0 , 0 , n122 );
and_AQFP n123_( clk_6 , splitterfromn116 , splitterfromn122 , 0 , 0 , n123 );
or_AQFP n124_( clk_6 , splitterfromn116 , splitterfromn122 , 0 , 0 , n124 );
and_AQFP n125_( clk_7 , n123 , n124 , 1 , 0 , n125 );
or_AQFP n126_( clk_1 , buf_splitterG31ton126n127_n126_2 , splitterfromn125 , 0 , 0 , n126 );
or_AQFP n127_( clk_5 , buf_splitterG23ton109n200_n127_4 , splitterG31ton126n127 , 0 , 0 , n127 );
and_AQFP n128_( clk_1 , buf_splitterfromG19_n128_5 , splitterfromn127 , 0 , 0 , n128 );
and_AQFP n129_( clk_3 , splitterfromn126 , splittern128ton129n295 , 0 , 0 , n129 );
or_AQFP n130_( clk_3 , splitterfromn126 , splittern128ton129n295 , 0 , 0 , n130 );
and_AQFP n131_( clk_4 , n129 , n130 , 1 , 0 , n131 );
and_AQFP n132_( clk_5 , n102 , n131 , 0 , 0 , n132 );
and_AQFP n133_( clk_6 , splitterfromG18 , splitterfromn88 , 0 , 1 , n133 );
or_AQFP n134_( clk_3 , splitterG11ton134n80 , splitterG15ton134n62 , 0 , 0 , n134 );
and_AQFP n135_( clk_3 , splitterG11ton134n80 , splitterG15ton134n62 , 0 , 0 , n135 );
and_AQFP n136_( clk_4 , n134 , n135 , 0 , 1 , n136 );
or_AQFP n137_( clk_8 , splitterfromn133 , splitterfromn136 , 0 , 0 , n137 );
and_AQFP n138_( clk_8 , splitterfromn133 , splitterfromn136 , 0 , 0 , n138 );
and_AQFP n139_( clk_1 , n137 , n138 , 0 , 1 , n139 );
and_AQFP n140_( clk_3 , splittern108ton114n141 , splitterfromn139 , 0 , 0 , n140 );
or_AQFP n141_( clk_3 , splittern108ton114n141 , splitterfromn139 , 0 , 0 , n141 );
and_AQFP n142_( clk_4 , n140 , n141 , 1 , 0 , n142 );
and_AQFP n143_( clk_3 , splitterG5ton143n40 , splitterG8ton143n43 , 0 , 1 , n143 );
and_AQFP n144_( clk_3 , splitterG5ton143n40 , splitterG8ton143n43 , 1 , 0 , n144 );
or_AQFP n145_( clk_4 , n143 , n144 , 0 , 0 , n145 );
and_AQFP n146_( clk_6 , buf_splitterG2ton146n46_n146_1 , splitterfromn145 , 0 , 1 , n146 );
and_AQFP n147_( clk_6 , buf_splitterG2ton146n46_n147_1 , splitterfromn145 , 1 , 0 , n147 );
or_AQFP n148_( clk_8 , n146 , n147 , 0 , 0 , n148 );
and_AQFP n149_( clk_6 , splitterfromn142 , splitterfromn148 , 1 , 0 , n149 );
and_AQFP n150_( clk_6 , splitterfromn142 , splitterfromn148 , 0 , 1 , n150 );
or_AQFP n151_( clk_7 , n149 , n150 , 0 , 0 , n151 );
and_AQFP n152_( clk_1 , buf_splitterG31ton152n201_n152_2 , splitterfromn151 , 1 , 0 , n152 );
and_AQFP n153_( clk_3 , splitterG27ton153n287 , splitterfromn152 , 0 , 0 , n153 );
or_AQFP n154_( clk_3 , splitterG27ton153n287 , splitterfromn152 , 0 , 0 , n154 );
and_AQFP n155_( clk_4 , n153 , n154 , 1 , 0 , n155 );
or_AQFP n156_( clk_4 , splitterG3ton156n46 , splitterG6ton156n37 , 0 , 0 , n156 );
and_AQFP n157_( clk_4 , splitterG3ton156n46 , splitterG6ton156n37 , 0 , 0 , n157 );
and_AQFP n158_( clk_6 , n156 , n157 , 0 , 1 , n158 );
and_AQFP n159_( clk_2 , splitterG8ton159n160 , splitterfromn158 , 0 , 0 , n159 );
or_AQFP n160_( clk_2 , splitterG8ton159n160 , splitterfromn158 , 0 , 0 , n160 );
and_AQFP n161_( clk_3 , n159 , n160 , 1 , 0 , n161 );
and_AQFP n162_( clk_7 , splitterfromG19 , splitterfromn109 , 0 , 1 , n162 );
and_AQFP n163_( clk_7 , splitterG12ton163n83 , splittern63ton163n65 , 0 , 0 , n163 );
or_AQFP n164_( clk_7 , splitterG12ton163n83 , splittern63ton163n65 , 0 , 0 , n164 );
and_AQFP n165_( clk_8 , n163 , n164 , 1 , 0 , n165 );
and_AQFP n166_( clk_2 , splitterfromn162 , splitterfromn165 , 0 , 1 , n166 );
and_AQFP n167_( clk_2 , splitterfromn162 , splitterfromn165 , 1 , 0 , n167 );
or_AQFP n168_( clk_3 , n166 , n167 , 0 , 0 , n168 );
or_AQFP n169_( clk_5 , splitterfromn161 , splitterfromn168 , 0 , 0 , n169 );
and_AQFP n170_( clk_5 , splitterfromn161 , splitterfromn168 , 0 , 0 , n170 );
and_AQFP n171_( clk_7 , n169 , n170 , 0 , 1 , n171 );
and_AQFP n172_( clk_1 , buf_splitterG31ton152n201_n172_1 , splitterfromn171 , 1 , 0 , n172 );
and_AQFP n173_( clk_3 , splitterG28ton173n291 , splitterfromn172 , 0 , 0 , n173 );
or_AQFP n174_( clk_3 , splitterG28ton173n291 , splitterfromn172 , 0 , 0 , n174 );
and_AQFP n175_( clk_4 , n173 , n174 , 1 , 0 , n175 );
or_AQFP n176_( clk_5 , n155 , n175 , 0 , 0 , n176 );
and_AQFP n177_( clk_6 , n132 , n176 , 0 , 1 , n177 );
and_AQFP n178_( clk_8 , buf_splitterfromG20_n178_6 , splitterfromn127 , 0 , 0 , n178 );
and_AQFP n179_( clk_5 , splitterfromG22 , buf_splitterG33ton109n88_n179_1 , 0 , 1 , n179 );
and_AQFP n180_( clk_5 , buf_splitterG14ton103n265_n180_1 , splitterG4ton180n181 , 1 , 0 , n180 );
and_AQFP n181_( clk_6 , splitterG14ton181n265 , splitterG4ton180n181 , 0 , 1 , n181 );
or_AQFP n182_( clk_7 , n180 , n181 , 0 , 0 , n182 );
and_AQFP n183_( clk_1 , splitterfromn179 , splitterfromn182 , 0 , 1 , n183 );
and_AQFP n184_( clk_1 , splitterfromn179 , splitterfromn182 , 1 , 0 , n184 );
or_AQFP n185_( clk_2 , n183 , n184 , 0 , 0 , n185 );
or_AQFP n186_( clk_4 , buf_splittern50ton186n52_n186_1 , splitterfromn185 , 0 , 0 , n186 );
and_AQFP n187_( clk_4 , buf_splittern50ton186n52_n187_1 , splitterfromn185 , 0 , 0 , n187 );
and_AQFP n188_( clk_5 , n186 , n187 , 0 , 1 , n188 );
or_AQFP n189_( clk_7 , buf_splittern87ton189n97_n189_1 , splitterfromn188 , 0 , 0 , n189 );
and_AQFP n190_( clk_7 , buf_splittern87ton189n97_n190_1 , splitterfromn188 , 0 , 0 , n190 );
and_AQFP n191_( clk_8 , n189 , n190 , 0 , 1 , n191 );
and_AQFP n192_( clk_2 , buf_splitterG31ton152n201_n192_2 , splitterfromn191 , 1 , 0 , n192 );
or_AQFP n193_( clk_4 , splitterG25ton193n281 , splittern192ton193n284 , 0 , 0 , n193 );
and_AQFP n194_( clk_4 , splitterG25ton193n281 , splittern192ton193n284 , 0 , 0 , n194 );
and_AQFP n195_( clk_5 , n193 , n194 , 0 , 1 , n195 );
and_AQFP n196_( clk_7 , splittern178ton196n269 , splittern195ton196n270 , 0 , 0 , n196 );
and_AQFP n197_( clk_8 , splittern177ton197n272 , n196 , 0 , 1 , n197 );
and_AQFP n198_( clk_2 , splitterfromn78 , splitterfromn197 , 1 , 0 , n198 );
or_AQFP n199_( clk_6 , buf_splitterfromG29_n199_1 , splitterG33ton199n273 , 0 , 0 , n199 );
and_AQFP n200_( clk_6 , buf_splitterG23ton109n200_n200_1 , buf_splitterG24ton200n88_n200_1 , 1 , 0 , n200 );
or_AQFP n201_( clk_6 , splitterG31ton152n201 , splitterfromn200 , 0 , 0 , n201 );
or_AQFP n202_( clk_8 , splitterfromn199 , splitterfromn201 , 0 , 0 , n202 );
or_AQFP n203_( clk_7 , splitterfromG32 , buf_splitterG33ton199n273_n203_1 , 0 , 0 , n203 );
or_AQFP n204_( clk_8 , buf_splitterfromn200_n204_1 , splittern203ton204n321 , 0 , 0 , n204 );
and_AQFP n205_( clk_3 , buf_n202_n205_1 , splitterfromn204 , 0 , 0 , n205 );
and_AQFP n206_( clk_4 , splitterfromn198 , buf_splitterfromn205_n206_4 , 0 , 1 , n206 );
or_AQFP n207_( clk_6 , buf_splitterG1ton207n91_n207_12 , splittern206ton207n302 , 0 , 0 , n207 );
and_AQFP n208_( clk_7 , buf_splitterG1ton207n91_n208_12 , splittern206ton208n210 , 0 , 0 , n208 );
and_AQFP n209_( clk_8 , n207 , n208 , 0 , 1 , n209 );
or_AQFP n210_( clk_8 , buf_splitterG2ton146n46_n210_14 , splittern206ton208n210 , 0 , 0 , n210 );
and_AQFP n211_( clk_8 , buf_splitterG2ton211n46_n211_14 , splittern206ton211n216 , 0 , 0 , n211 );
and_AQFP n212_( clk_2 , n210 , n211 , 0 , 1 , n212 );
or_AQFP n213_( clk_8 , buf_splitterG3ton156n46_n213_15 , splittern206ton211n216 , 0 , 0 , n213 );
and_AQFP n214_( clk_7 , buf_splitterG3ton214n46_n214_13 , splittern206ton211n216 , 0 , 0 , n214 );
and_AQFP n215_( clk_2 , n213 , buf_n214_n215_1 , 0 , 1 , n215 );
or_AQFP n216_( clk_8 , buf_splitterG4ton216n43_n216_13 , splittern206ton211n216 , 0 , 0 , n216 );
and_AQFP n217_( clk_7 , buf_splitterG4ton216n43_n217_12 , splittern206ton217n302 , 0 , 0 , n217 );
and_AQFP n218_( clk_1 , n216 , n217 , 0 , 1 , n218 );
or_AQFP n219_( clk_5 , splitterfromG30 , splitterG33ton199n273 , 0 , 0 , n219 );
or_AQFP n220_( clk_8 , splitterfromn201 , splitterfromn219 , 0 , 0 , n220 );
and_AQFP n221_( clk_2 , splitterfromn204 , n220 , 0 , 0 , n221 );
and_AQFP n222_( clk_4 , splitterfromn198 , buf_splittern221ton222n254_n222_2 , 0 , 1 , n222 );
or_AQFP n223_( clk_6 , buf_splitterG10ton120n62_n223_13 , splittern222ton223n314 , 0 , 0 , n223 );
and_AQFP n224_( clk_6 , buf_splitterG10ton224n62_n224_13 , splittern222ton223n314 , 0 , 0 , n224 );
and_AQFP n225_( clk_8 , n223 , n224 , 0 , 1 , n225 );
or_AQFP n226_( clk_7 , buf_splitterG15ton134n62_n226_14 , splittern222ton226n229 , 0 , 0 , n226 );
and_AQFP n227_( clk_8 , buf_splitterG15ton227n62_n227_14 , splittern222ton226n229 , 0 , 0 , n227 );
and_AQFP n228_( clk_2 , buf_n226_n228_1 , n227 , 0 , 1 , n228 );
or_AQFP n229_( clk_7 , buf_splitterG16ton106n65_n229_13 , splittern222ton226n229 , 0 , 0 , n229 );
and_AQFP n230_( clk_8 , buf_splitterG16ton230n65_n230_12 , splittern222ton230n314 , 0 , 0 , n230 );
and_AQFP n231_( clk_1 , n229 , n230 , 0 , 1 , n231 );
and_AQFP n232_( clk_7 , splittern178ton196n269 , splittern195ton196n270 , 0 , 1 , n232 );
and_AQFP n233_( clk_8 , splittern177ton197n272 , n232 , 0 , 0 , n233 );
and_AQFP n234_( clk_2 , splitterfromn78 , n233 , 1 , 0 , n234 );
and_AQFP n235_( clk_4 , buf_splitterfromn205_n235_6 , splitterfromn234 , 1 , 0 , n235 );
or_AQFP n236_( clk_6 , buf_splitterG5ton143n40_n236_13 , splittern235ton236n246 , 0 , 0 , n236 );
and_AQFP n237_( clk_6 , buf_splitterG5ton237n40_n237_11 , splittern235ton236n246 , 0 , 0 , n237 );
and_AQFP n238_( clk_8 , n236 , n237 , 0 , 1 , n238 );
or_AQFP n239_( clk_8 , buf_splitterG6ton156n37_n239_14 , splittern235ton239n240 , 0 , 0 , n239 );
and_AQFP n240_( clk_7 , buf_splitterG6ton240n37_n240_13 , splittern235ton239n240 , 0 , 0 , n240 );
and_AQFP n241_( clk_1 , n239 , n240 , 0 , 1 , n241 );
or_AQFP n242_( clk_8 , buf_splitterG7ton117n37_n242_14 , splittern235ton242n246 , 0 , 0 , n242 );
and_AQFP n243_( clk_7 , buf_splitterG7ton243n37_n243_15 , splittern235ton242n246 , 0 , 0 , n243 );
and_AQFP n244_( clk_2 , n242 , buf_n243_n244_1 , 0 , 1 , n244 );
or_AQFP n245_( clk_7 , buf_splitterG8ton245n43_n245_12 , splittern235ton242n246 , 0 , 0 , n245 );
and_AQFP n246_( clk_7 , buf_splitterG8ton245n43_n246_12 , splittern235ton242n246 , 0 , 0 , n246 );
and_AQFP n247_( clk_8 , n245 , n246 , 0 , 1 , n247 );
and_AQFP n248_( clk_4 , buf_splittern221ton222n254_n248_2 , splitterfromn234 , 1 , 0 , n248 );
and_AQFP n249_( clk_6 , buf_splitterG9ton103n59_n249_13 , splitterfromn248 , 0 , 1 , n249 );
and_AQFP n250_( clk_6 , buf_splitterG9ton250n59_n250_11 , splitterfromn248 , 1 , 0 , n250 );
or_AQFP n251_( clk_7 , n249 , n250 , 0 , 0 , n251 );
and_AQFP n252_( clk_2 , buf_splittern35ton252n78_n252_2 , splitterfromn197 , 0 , 0 , n252 );
and_AQFP n253_( clk_3 , buf_splittern77ton253n78_n253_1 , n252 , 0 , 0 , n253 );
and_AQFP n254_( clk_4 , buf_splittern221ton222n254_n254_2 , n253 , 1 , 0 , n254 );
or_AQFP n255_( clk_6 , buf_splitterG11ton134n80_n255_13 , splittern254ton255n265 , 0 , 0 , n255 );
and_AQFP n256_( clk_6 , buf_splitterG11ton256n80_n256_13 , splittern254ton255n265 , 0 , 0 , n256 );
and_AQFP n257_( clk_8 , n255 , n256 , 0 , 1 , n257 );
or_AQFP n258_( clk_7 , buf_splitterG12ton163n83_n258_13 , splittern254ton258n259 , 0 , 0 , n258 );
and_AQFP n259_( clk_7 , buf_splitterG12ton259n83_n259_12 , splittern254ton258n259 , 0 , 0 , n259 );
and_AQFP n260_( clk_8 , n258 , n259 , 0 , 1 , n260 );
or_AQFP n261_( clk_8 , buf_splitterG13ton111n80_n261_15 , splittern254ton261n265 , 0 , 0 , n261 );
and_AQFP n262_( clk_8 , buf_splitterG13ton262n80_n262_14 , splittern254ton261n265 , 0 , 0 , n262 );
and_AQFP n263_( clk_2 , n261 , n262 , 0 , 1 , n263 );
or_AQFP n264_( clk_7 , buf_splitterG14ton181n265_n264_13 , splittern254ton261n265 , 0 , 0 , n264 );
and_AQFP n265_( clk_7 , buf_splitterG14ton181n265_n265_13 , splittern254ton261n265 , 0 , 0 , n265 );
and_AQFP n266_( clk_8 , n264 , n265 , 0 , 1 , n266 );
or_AQFP n267_( clk_7 , splittern206ton217n302 , splittern222ton230n314 , 0 , 0 , n267 );
and_AQFP n268_( clk_1 , buf_splitterfromG32_n268_14 , splittern267ton268n320 , 0 , 0 , n268 );
or_AQFP n269_( clk_6 , splittern35ton252n78 , splittern178ton196n269 , 0 , 0 , n269 );
or_AQFP n270_( clk_7 , splittern195ton196n270 , n269 , 0 , 0 , n270 );
and_AQFP n271_( clk_8 , splittern77ton253n78 , n270 , 0 , 1 , n271 );
and_AQFP n272_( clk_2 , buf_splittern177ton197n272_n272_1 , n271 , 0 , 0 , n272 );
or_AQFP n273_( clk_4 , buf_splitterG33ton199n273_n273_11 , n272 , 0 , 0 , n273 );
or_AQFP n274_( clk_2 , n268 , buf_n273_n274_3 , 0 , 0 , n274 );
and_AQFP n275_( clk_1 , buf_splittern74ton275n76_n275_8 , splittern267ton268n320 , 0 , 0 , n275 );
and_AQFP n276_( clk_3 , buf_splitterG31ton276n291_n276_8 , splitterfromn275 , 1 , 0 , n276 );
and_AQFP n277_( clk_4 , buf_splitterfromn72_n277_9 , n276 , 0 , 1 , n277 );
and_AQFP n278_( clk_3 , buf_splittern73ton278n76_n278_7 , splitterfromn275 , 1 , 0 , n278 );
and_AQFP n279_( clk_4 , buf_splittern203ton204n321_n279_13 , n278 , 0 , 1 , n279 );
and_AQFP n280_( clk_5 , n277 , n279 , 1 , 0 , n280 );
and_AQFP n281_( clk_1 , buf_splitterG25ton193n281_n281_9 , splittern267ton268n320 , 0 , 0 , n281 );
and_AQFP n282_( clk_3 , buf_splitterG31ton276n291_n282_8 , splitterfromn281 , 1 , 0 , n282 );
or_AQFP n283_( clk_4 , buf_splitterfromn191_n283_10 , n282 , 0 , 0 , n283 );
and_AQFP n284_( clk_3 , buf_splittern192ton193n284_n284_7 , splitterfromn281 , 0 , 0 , n284 );
and_AQFP n285_( clk_4 , buf_splittern203ton204n321_n285_14 , n284 , 0 , 1 , n285 );
and_AQFP n286_( clk_5 , n283 , n285 , 0 , 0 , n286 );
and_AQFP n287_( clk_4 , buf_splitterG27ton153n287_n287_1 , splitterG31ton276n291 , 0 , 1 , n287 );
and_AQFP n288_( clk_3 , splittern267ton288n320 , buf_n287_n288_7 , 0 , 0 , n288 );
and_AQFP n289_( clk_4 , buf_splitterfromn151_n289_9 , n288 , 0 , 1 , n289 );
and_AQFP n290_( clk_5 , buf_splittern203ton290n321_n290_1 , n289 , 0 , 1 , n290 );
and_AQFP n291_( clk_5 , buf_splitterG28ton173n291_n291_1 , splitterG31ton276n291 , 0 , 1 , n291 );
and_AQFP n292_( clk_2 , splittern267ton288n320 , buf_n291_n292_6 , 0 , 0 , n292 );
and_AQFP n293_( clk_3 , buf_splitterfromn171_n293_9 , n292 , 0 , 1 , n293 );
and_AQFP n294_( clk_4 , buf_splittern203ton290n321_n294_1 , n293 , 0 , 1 , n294 );
and_AQFP n295_( clk_6 , buf_splitterG31ton295n99_n295_5 , buf_splittern128ton129n295_n295_1 , 1 , 0 , n295 );
and_AQFP n296_( clk_2 , splittern267ton288n320 , buf_n295_n296_5 , 0 , 0 , n296 );
or_AQFP n297_( clk_3 , buf_splitterfromn125_n297_10 , n296 , 0 , 0 , n297 );
and_AQFP n298_( clk_4 , splittern203ton290n321 , n297 , 0 , 0 , n298 );
and_AQFP n299_( clk_8 , splittern56ton299n71 , splitterfromn199 , 0 , 0 , n299 );
and_AQFP n300_( clk_5 , splitterfromG21 , splitterfromG29 , 0 , 0 , n300 );
or_AQFP n301_( clk_7 , splittern206ton217n302 , buf_splitterfromn300_n301_9 , 0 , 0 , n301 );
and_AQFP n302_( clk_7 , splittern206ton217n302 , buf_splitterfromn300_n302_10 , 0 , 0 , n302 );
and_AQFP n303_( clk_8 , n301 , n302 , 0 , 1 , n303 );
or_AQFP n304_( clk_1 , buf_splitterG33ton304n88_n304_14 , n303 , 0 , 0 , n304 );
and_AQFP n305_( clk_3 , buf_splitterfromn299_n305_8 , splitterfromn304 , 0 , 0 , n305 );
or_AQFP n306_( clk_3 , buf_splitterfromn299_n306_8 , splitterfromn304 , 0 , 0 , n306 );
and_AQFP n307_( clk_5 , n305 , n306 , 1 , 0 , n307 );
or_AQFP n308_( clk_5 , splittern87ton189n97 , buf_splittern105ton106n309_n308_3 , 0 , 0 , n308 );
and_AQFP n309_( clk_6 , splittern87ton309n97 , buf_splittern105ton106n309_n309_4 , 0 , 0 , n309 );
and_AQFP n310_( clk_2 , buf_splitterfromn219_n310_1 , buf_n309_n310_1 , 0 , 1 , n310 );
and_AQFP n311_( clk_3 , buf_n308_n311_2 , n310 , 0 , 0 , n311 );
and_AQFP n312_( clk_6 , splitterfromG22 , buf_splitterfromG30_n312_1 , 0 , 0 , n312 );
or_AQFP n313_( clk_7 , splittern222ton230n314 , buf_splitterfromn312_n313_10 , 0 , 0 , n313 );
and_AQFP n314_( clk_7 , splittern222ton230n314 , buf_splitterfromn312_n314_12 , 0 , 0 , n314 );
and_AQFP n315_( clk_8 , n313 , n314 , 0 , 1 , n315 );
or_AQFP n316_( clk_1 , buf_splitterG33ton304n88_n316_16 , n315 , 0 , 0 , n316 );
and_AQFP n317_( clk_3 , buf_splitterfromn311_n317_3 , splitterfromn316 , 0 , 1 , n317 );
and_AQFP n318_( clk_3 , buf_splitterfromn311_n318_4 , splitterfromn316 , 1 , 0 , n318 );
or_AQFP n319_( clk_5 , n317 , n318 , 0 , 0 , n319 );
and_AQFP n320_( clk_2 , buf_splitterG26ton100n320_n320_8 , splittern267ton288n320 , 0 , 0 , n320 );
and_AQFP n321_( clk_3 , buf_splitterfromn98_n321_10 , splittern203ton290n321 , 1 , 0 , n321 );
and_AQFP n322_( clk_4 , n320 , n321 , 1 , 0 , n322 );
PO_AQFP G1884_( clk_6 , buf_n209_G1884_2 , 1 , G1884 );
PO_AQFP G1885_( clk_6 , buf_n212_G1885_1 , 1 , G1885 );
PO_AQFP G1886_( clk_6 , buf_n215_G1886_1 , 1 , G1886 );
PO_AQFP G1887_( clk_6 , buf_n218_G1887_2 , 1 , G1887 );
PO_AQFP G1888_( clk_6 , buf_n225_G1888_4 , 1 , G1888 );
PO_AQFP G1889_( clk_6 , buf_n228_G1889_1 , 1 , G1889 );
PO_AQFP G1890_( clk_6 , buf_n231_G1890_2 , 1 , G1890 );
PO_AQFP G1891_( clk_6 , buf_n238_G1891_2 , 1 , G1891 );
PO_AQFP G1892_( clk_6 , buf_n241_G1892_2 , 1 , G1892 );
PO_AQFP G1893_( clk_6 , buf_n244_G1893_1 , 1 , G1893 );
PO_AQFP G1894_( clk_6 , buf_n247_G1894_3 , 1 , G1894 );
PO_AQFP G1895_( clk_6 , buf_n251_G1895_5 , 1 , G1895 );
PO_AQFP G1896_( clk_6 , buf_n257_G1896_2 , 1 , G1896 );
PO_AQFP G1897_( clk_6 , buf_n260_G1897_4 , 1 , G1897 );
PO_AQFP G1898_( clk_6 , buf_n263_G1898_1 , 1 , G1898 );
PO_AQFP G1899_( clk_6 , buf_n266_G1899_3 , 1 , G1899 );
PO_AQFP G1900_( clk_6 , buf_n274_G1900_1 , 0 , G1900 );
PO_AQFP G1901_( clk_6 , n280 , 0 , G1901 );
PO_AQFP G1902_( clk_6 , n286 , 0 , G1902 );
PO_AQFP G1903_( clk_6 , n290 , 0 , G1903 );
PO_AQFP G1904_( clk_6 , n294 , 0 , G1904 );
PO_AQFP G1905_( clk_6 , n298 , 0 , G1905 );
PO_AQFP G1906_( clk_6 , n307 , 1 , G1906 );
PO_AQFP G1907_( clk_6 , n319 , 1 , G1907 );
PO_AQFP G1908_( clk_6 , n322 , 0 , G1908 );
buf_AQFP buf_G1_splitterG1ton207n91_1_( clk_2 , G1 , 0 , buf_G1_splitterG1ton207n91_1 );
buf_AQFP buf_G1_splitterG1ton207n91_2_( clk_3 , buf_G1_splitterG1ton207n91_1 , 0 , buf_G1_splitterG1ton207n91_2 );
buf_AQFP buf_G12_splitterG12ton163n83_1_( clk_3 , G12 , 0 , buf_G12_splitterG12ton163n83_1 );
buf_AQFP buf_G16_splitterG16ton106n65_1_( clk_2 , G16 , 0 , buf_G16_splitterG16ton106n65_1 );
buf_AQFP buf_G16_splitterG16ton106n65_2_( clk_3 , buf_G16_splitterG16ton106n65_1 , 0 , buf_G16_splitterG16ton106n65_2 );
buf_AQFP buf_G17_splitterfromG17_1_( clk_2 , G17 , 0 , buf_G17_splitterfromG17_1 );
buf_AQFP buf_G18_splitterfromG18_1_( clk_3 , G18 , 0 , buf_G18_splitterfromG18_1 );
buf_AQFP buf_G19_splitterfromG19_1_( clk_2 , G19 , 0 , buf_G19_splitterfromG19_1 );
buf_AQFP buf_G19_splitterfromG19_2_( clk_4 , buf_G19_splitterfromG19_1 , 0 , buf_G19_splitterfromG19_2 );
buf_AQFP buf_G20_splitterfromG20_1_( clk_2 , G20 , 0 , buf_G20_splitterfromG20_1 );
buf_AQFP buf_G22_splitterfromG22_1_( clk_2 , G22 , 0 , buf_G22_splitterfromG22_1 );
buf_AQFP buf_G24_splitterG24ton200n88_1_( clk_2 , G24 , 0 , buf_G24_splitterG24ton200n88_1 );
buf_AQFP buf_G25_splitterG25ton193n281_1_( clk_3 , G25 , 0 , buf_G25_splitterG25ton193n281_1 );
buf_AQFP buf_G25_splitterG25ton193n281_2_( clk_5 , buf_G25_splitterG25ton193n281_1 , 0 , buf_G25_splitterG25ton193n281_2 );
buf_AQFP buf_G25_splitterG25ton193n281_3_( clk_7 , buf_G25_splitterG25ton193n281_2 , 0 , buf_G25_splitterG25ton193n281_3 );
buf_AQFP buf_G25_splitterG25ton193n281_4_( clk_1 , buf_G25_splitterG25ton193n281_3 , 0 , buf_G25_splitterG25ton193n281_4 );
buf_AQFP buf_G25_splitterG25ton193n281_5_( clk_3 , buf_G25_splitterG25ton193n281_4 , 0 , buf_G25_splitterG25ton193n281_5 );
buf_AQFP buf_G25_splitterG25ton193n281_6_( clk_5 , buf_G25_splitterG25ton193n281_5 , 0 , buf_G25_splitterG25ton193n281_6 );
buf_AQFP buf_G25_splitterG25ton193n281_7_( clk_6 , buf_G25_splitterG25ton193n281_6 , 0 , buf_G25_splitterG25ton193n281_7 );
buf_AQFP buf_G25_splitterG25ton193n281_8_( clk_8 , buf_G25_splitterG25ton193n281_7 , 0 , buf_G25_splitterG25ton193n281_8 );
buf_AQFP buf_G25_splitterG25ton193n281_9_( clk_1 , buf_G25_splitterG25ton193n281_8 , 0 , buf_G25_splitterG25ton193n281_9 );
buf_AQFP buf_G26_splitterG26ton100n320_1_( clk_3 , G26 , 0 , buf_G26_splitterG26ton100n320_1 );
buf_AQFP buf_G26_splitterG26ton100n320_2_( clk_5 , buf_G26_splitterG26ton100n320_1 , 0 , buf_G26_splitterG26ton100n320_2 );
buf_AQFP buf_G26_splitterG26ton100n320_3_( clk_7 , buf_G26_splitterG26ton100n320_2 , 0 , buf_G26_splitterG26ton100n320_3 );
buf_AQFP buf_G26_splitterG26ton100n320_4_( clk_1 , buf_G26_splitterG26ton100n320_3 , 0 , buf_G26_splitterG26ton100n320_4 );
buf_AQFP buf_G26_splitterG26ton100n320_5_( clk_3 , buf_G26_splitterG26ton100n320_4 , 0 , buf_G26_splitterG26ton100n320_5 );
buf_AQFP buf_G26_splitterG26ton100n320_6_( clk_5 , buf_G26_splitterG26ton100n320_5 , 0 , buf_G26_splitterG26ton100n320_6 );
buf_AQFP buf_G26_splitterG26ton100n320_7_( clk_7 , buf_G26_splitterG26ton100n320_6 , 0 , buf_G26_splitterG26ton100n320_7 );
buf_AQFP buf_G27_splitterG27ton153n287_1_( clk_3 , G27 , 0 , buf_G27_splitterG27ton153n287_1 );
buf_AQFP buf_G27_splitterG27ton153n287_2_( clk_5 , buf_G27_splitterG27ton153n287_1 , 0 , buf_G27_splitterG27ton153n287_2 );
buf_AQFP buf_G27_splitterG27ton153n287_3_( clk_7 , buf_G27_splitterG27ton153n287_2 , 0 , buf_G27_splitterG27ton153n287_3 );
buf_AQFP buf_G27_splitterG27ton153n287_4_( clk_1 , buf_G27_splitterG27ton153n287_3 , 0 , buf_G27_splitterG27ton153n287_4 );
buf_AQFP buf_G27_splitterG27ton153n287_5_( clk_3 , buf_G27_splitterG27ton153n287_4 , 0 , buf_G27_splitterG27ton153n287_5 );
buf_AQFP buf_G27_splitterG27ton153n287_6_( clk_5 , buf_G27_splitterG27ton153n287_5 , 0 , buf_G27_splitterG27ton153n287_6 );
buf_AQFP buf_G27_splitterG27ton153n287_7_( clk_7 , buf_G27_splitterG27ton153n287_6 , 0 , buf_G27_splitterG27ton153n287_7 );
buf_AQFP buf_G28_splitterG28ton173n291_1_( clk_2 , G28 , 0 , buf_G28_splitterG28ton173n291_1 );
buf_AQFP buf_G28_splitterG28ton173n291_2_( clk_3 , buf_G28_splitterG28ton173n291_1 , 0 , buf_G28_splitterG28ton173n291_2 );
buf_AQFP buf_G28_splitterG28ton173n291_3_( clk_5 , buf_G28_splitterG28ton173n291_2 , 0 , buf_G28_splitterG28ton173n291_3 );
buf_AQFP buf_G28_splitterG28ton173n291_4_( clk_7 , buf_G28_splitterG28ton173n291_3 , 0 , buf_G28_splitterG28ton173n291_4 );
buf_AQFP buf_G28_splitterG28ton173n291_5_( clk_1 , buf_G28_splitterG28ton173n291_4 , 0 , buf_G28_splitterG28ton173n291_5 );
buf_AQFP buf_G28_splitterG28ton173n291_6_( clk_3 , buf_G28_splitterG28ton173n291_5 , 0 , buf_G28_splitterG28ton173n291_6 );
buf_AQFP buf_G28_splitterG28ton173n291_7_( clk_5 , buf_G28_splitterG28ton173n291_6 , 0 , buf_G28_splitterG28ton173n291_7 );
buf_AQFP buf_G28_splitterG28ton173n291_8_( clk_7 , buf_G28_splitterG28ton173n291_7 , 0 , buf_G28_splitterG28ton173n291_8 );
buf_AQFP buf_G29_splitterfromG29_1_( clk_2 , G29 , 0 , buf_G29_splitterfromG29_1 );
buf_AQFP buf_G30_splitterfromG30_1_( clk_2 , G30 , 0 , buf_G30_splitterfromG30_1 );
buf_AQFP buf_G32_splitterfromG32_1_( clk_2 , G32 , 0 , buf_G32_splitterfromG32_1 );
buf_AQFP buf_G32_splitterfromG32_2_( clk_3 , buf_G32_splitterfromG32_1 , 0 , buf_G32_splitterfromG32_2 );
buf_AQFP buf_G32_splitterfromG32_3_( clk_5 , buf_G32_splitterfromG32_2 , 0 , buf_G32_splitterfromG32_3 );
buf_AQFP buf_n35_splittern35ton252n78_1_( clk_6 , n35 , 0 , buf_n35_splittern35ton252n78_1 );
buf_AQFP buf_n35_splittern35ton252n78_2_( clk_8 , buf_n35_splittern35ton252n78_1 , 0 , buf_n35_splittern35ton252n78_2 );
buf_AQFP buf_n35_splittern35ton252n78_3_( clk_2 , buf_n35_splittern35ton252n78_2 , 0 , buf_n35_splittern35ton252n78_3 );
buf_AQFP buf_n57_splitterfromn57_1_( clk_6 , n57 , 0 , buf_n57_splitterfromn57_1 );
buf_AQFP buf_n74_splittern74ton275n76_1_( clk_1 , n74 , 0 , buf_n74_splittern74ton275n76_1 );
buf_AQFP buf_n122_splitterfromn122_1_( clk_2 , n122 , 0 , buf_n122_splitterfromn122_1 );
buf_AQFP buf_n148_splitterfromn148_1_( clk_1 , n148 , 0 , buf_n148_splitterfromn148_1 );
buf_AQFP buf_n148_splitterfromn148_2_( clk_2 , buf_n148_splitterfromn148_1 , 0 , buf_n148_splitterfromn148_2 );
buf_AQFP buf_n178_splittern178ton196n269_1_( clk_1 , n178 , 0 , buf_n178_splittern178ton196n269_1 );
buf_AQFP buf_n178_splittern178ton196n269_2_( clk_3 , buf_n178_splittern178ton196n269_1 , 0 , buf_n178_splittern178ton196n269_2 );
buf_AQFP buf_n199_splitterfromn199_1_( clk_8 , n199 , 0 , buf_n199_splitterfromn199_1 );
buf_AQFP buf_n199_splitterfromn199_2_( clk_2 , buf_n199_splitterfromn199_1 , 0 , buf_n199_splitterfromn199_2 );
buf_AQFP buf_n199_splitterfromn199_3_( clk_4 , buf_n199_splitterfromn199_2 , 0 , buf_n199_splitterfromn199_3 );
buf_AQFP buf_n200_splitterfromn200_1_( clk_8 , n200 , 0 , buf_n200_splitterfromn200_1 );
buf_AQFP buf_n200_splitterfromn200_2_( clk_2 , buf_n200_splitterfromn200_1 , 0 , buf_n200_splitterfromn200_2 );
buf_AQFP buf_n202_n205_1_( clk_1 , n202 , 0 , buf_n202_n205_1 );
buf_AQFP buf_n203_splittern203ton204n321_1_( clk_1 , n203 , 0 , buf_n203_splittern203ton204n321_1 );
buf_AQFP buf_n203_splittern203ton204n321_2_( clk_3 , buf_n203_splittern203ton204n321_1 , 0 , buf_n203_splittern203ton204n321_2 );
buf_AQFP buf_n203_splittern203ton204n321_3_( clk_4 , buf_n203_splittern203ton204n321_2 , 0 , buf_n203_splittern203ton204n321_3 );
buf_AQFP buf_n209_G1884_1_( clk_2 , n209 , 0 , buf_n209_G1884_1 );
buf_AQFP buf_n209_G1884_2_( clk_4 , buf_n209_G1884_1 , 0 , buf_n209_G1884_2 );
buf_AQFP buf_n212_G1885_1_( clk_4 , n212 , 0 , buf_n212_G1885_1 );
buf_AQFP buf_n214_n215_1_( clk_1 , n214 , 0 , buf_n214_n215_1 );
buf_AQFP buf_n215_G1886_1_( clk_4 , n215 , 0 , buf_n215_G1886_1 );
buf_AQFP buf_n218_G1887_1_( clk_3 , n218 , 0 , buf_n218_G1887_1 );
buf_AQFP buf_n218_G1887_2_( clk_5 , buf_n218_G1887_1 , 0 , buf_n218_G1887_2 );
buf_AQFP buf_n219_splitterfromn219_1_( clk_6 , n219 , 0 , buf_n219_splitterfromn219_1 );
buf_AQFP buf_n219_splitterfromn219_2_( clk_8 , buf_n219_splitterfromn219_1 , 0 , buf_n219_splitterfromn219_2 );
buf_AQFP buf_n219_splitterfromn219_3_( clk_1 , buf_n219_splitterfromn219_2 , 0 , buf_n219_splitterfromn219_3 );
buf_AQFP buf_n219_splitterfromn219_4_( clk_3 , buf_n219_splitterfromn219_3 , 0 , buf_n219_splitterfromn219_4 );
buf_AQFP buf_n219_splitterfromn219_5_( clk_5 , buf_n219_splitterfromn219_4 , 0 , buf_n219_splitterfromn219_5 );
buf_AQFP buf_n221_splittern221ton222n254_1_( clk_4 , n221 , 0 , buf_n221_splittern221ton222n254_1 );
buf_AQFP buf_n221_splittern221ton222n254_2_( clk_5 , buf_n221_splittern221ton222n254_1 , 0 , buf_n221_splittern221ton222n254_2 );
buf_AQFP buf_n225_G1888_1_( clk_1 , n225 , 0 , buf_n225_G1888_1 );
buf_AQFP buf_n225_G1888_2_( clk_2 , buf_n225_G1888_1 , 0 , buf_n225_G1888_2 );
buf_AQFP buf_n225_G1888_3_( clk_3 , buf_n225_G1888_2 , 0 , buf_n225_G1888_3 );
buf_AQFP buf_n225_G1888_4_( clk_4 , buf_n225_G1888_3 , 0 , buf_n225_G1888_4 );
buf_AQFP buf_n226_n228_1_( clk_1 , n226 , 0 , buf_n226_n228_1 );
buf_AQFP buf_n228_G1889_1_( clk_4 , n228 , 0 , buf_n228_G1889_1 );
buf_AQFP buf_n231_G1890_1_( clk_3 , n231 , 0 , buf_n231_G1890_1 );
buf_AQFP buf_n231_G1890_2_( clk_5 , buf_n231_G1890_1 , 0 , buf_n231_G1890_2 );
buf_AQFP buf_n238_G1891_1_( clk_2 , n238 , 0 , buf_n238_G1891_1 );
buf_AQFP buf_n238_G1891_2_( clk_4 , buf_n238_G1891_1 , 0 , buf_n238_G1891_2 );
buf_AQFP buf_n241_G1892_1_( clk_3 , n241 , 0 , buf_n241_G1892_1 );
buf_AQFP buf_n241_G1892_2_( clk_5 , buf_n241_G1892_1 , 0 , buf_n241_G1892_2 );
buf_AQFP buf_n243_n244_1_( clk_8 , n243 , 0 , buf_n243_n244_1 );
buf_AQFP buf_n244_G1893_1_( clk_4 , n244 , 0 , buf_n244_G1893_1 );
buf_AQFP buf_n247_G1894_1_( clk_1 , n247 , 0 , buf_n247_G1894_1 );
buf_AQFP buf_n247_G1894_2_( clk_3 , buf_n247_G1894_1 , 0 , buf_n247_G1894_2 );
buf_AQFP buf_n247_G1894_3_( clk_4 , buf_n247_G1894_2 , 0 , buf_n247_G1894_3 );
buf_AQFP buf_n251_G1895_1_( clk_8 , n251 , 0 , buf_n251_G1895_1 );
buf_AQFP buf_n251_G1895_2_( clk_1 , buf_n251_G1895_1 , 0 , buf_n251_G1895_2 );
buf_AQFP buf_n251_G1895_3_( clk_2 , buf_n251_G1895_2 , 0 , buf_n251_G1895_3 );
buf_AQFP buf_n251_G1895_4_( clk_3 , buf_n251_G1895_3 , 0 , buf_n251_G1895_4 );
buf_AQFP buf_n251_G1895_5_( clk_5 , buf_n251_G1895_4 , 0 , buf_n251_G1895_5 );
buf_AQFP buf_n257_G1896_1_( clk_2 , n257 , 0 , buf_n257_G1896_1 );
buf_AQFP buf_n257_G1896_2_( clk_4 , buf_n257_G1896_1 , 0 , buf_n257_G1896_2 );
buf_AQFP buf_n260_G1897_1_( clk_1 , n260 , 0 , buf_n260_G1897_1 );
buf_AQFP buf_n260_G1897_2_( clk_2 , buf_n260_G1897_1 , 0 , buf_n260_G1897_2 );
buf_AQFP buf_n260_G1897_3_( clk_3 , buf_n260_G1897_2 , 0 , buf_n260_G1897_3 );
buf_AQFP buf_n260_G1897_4_( clk_5 , buf_n260_G1897_3 , 0 , buf_n260_G1897_4 );
buf_AQFP buf_n263_G1898_1_( clk_4 , n263 , 0 , buf_n263_G1898_1 );
buf_AQFP buf_n266_G1899_1_( clk_1 , n266 , 0 , buf_n266_G1899_1 );
buf_AQFP buf_n266_G1899_2_( clk_2 , buf_n266_G1899_1 , 0 , buf_n266_G1899_2 );
buf_AQFP buf_n266_G1899_3_( clk_4 , buf_n266_G1899_2 , 0 , buf_n266_G1899_3 );
buf_AQFP buf_n273_n274_1_( clk_5 , n273 , 0 , buf_n273_n274_1 );
buf_AQFP buf_n273_n274_2_( clk_6 , buf_n273_n274_1 , 0 , buf_n273_n274_2 );
buf_AQFP buf_n273_n274_3_( clk_8 , buf_n273_n274_2 , 0 , buf_n273_n274_3 );
buf_AQFP buf_n274_G1900_1_( clk_4 , n274 , 0 , buf_n274_G1900_1 );
buf_AQFP buf_n287_n288_1_( clk_6 , n287 , 0 , buf_n287_n288_1 );
buf_AQFP buf_n287_n288_2_( clk_8 , buf_n287_n288_1 , 0 , buf_n287_n288_2 );
buf_AQFP buf_n287_n288_3_( clk_2 , buf_n287_n288_2 , 0 , buf_n287_n288_3 );
buf_AQFP buf_n287_n288_4_( clk_3 , buf_n287_n288_3 , 0 , buf_n287_n288_4 );
buf_AQFP buf_n287_n288_5_( clk_5 , buf_n287_n288_4 , 0 , buf_n287_n288_5 );
buf_AQFP buf_n287_n288_6_( clk_7 , buf_n287_n288_5 , 0 , buf_n287_n288_6 );
buf_AQFP buf_n287_n288_7_( clk_1 , buf_n287_n288_6 , 0 , buf_n287_n288_7 );
buf_AQFP buf_n291_n292_1_( clk_6 , n291 , 0 , buf_n291_n292_1 );
buf_AQFP buf_n291_n292_2_( clk_8 , buf_n291_n292_1 , 0 , buf_n291_n292_2 );
buf_AQFP buf_n291_n292_3_( clk_2 , buf_n291_n292_2 , 0 , buf_n291_n292_3 );
buf_AQFP buf_n291_n292_4_( clk_4 , buf_n291_n292_3 , 0 , buf_n291_n292_4 );
buf_AQFP buf_n291_n292_5_( clk_6 , buf_n291_n292_4 , 0 , buf_n291_n292_5 );
buf_AQFP buf_n291_n292_6_( clk_8 , buf_n291_n292_5 , 0 , buf_n291_n292_6 );
buf_AQFP buf_n295_n296_1_( clk_8 , n295 , 0 , buf_n295_n296_1 );
buf_AQFP buf_n295_n296_2_( clk_2 , buf_n295_n296_1 , 0 , buf_n295_n296_2 );
buf_AQFP buf_n295_n296_3_( clk_4 , buf_n295_n296_2 , 0 , buf_n295_n296_3 );
buf_AQFP buf_n295_n296_4_( clk_6 , buf_n295_n296_3 , 0 , buf_n295_n296_4 );
buf_AQFP buf_n295_n296_5_( clk_8 , buf_n295_n296_4 , 0 , buf_n295_n296_5 );
buf_AQFP buf_n300_splitterfromn300_1_( clk_6 , n300 , 0 , buf_n300_splitterfromn300_1 );
buf_AQFP buf_n300_splitterfromn300_2_( clk_8 , buf_n300_splitterfromn300_1 , 0 , buf_n300_splitterfromn300_2 );
buf_AQFP buf_n300_splitterfromn300_3_( clk_1 , buf_n300_splitterfromn300_2 , 0 , buf_n300_splitterfromn300_3 );
buf_AQFP buf_n300_splitterfromn300_4_( clk_2 , buf_n300_splitterfromn300_3 , 0 , buf_n300_splitterfromn300_4 );
buf_AQFP buf_n300_splitterfromn300_5_( clk_4 , buf_n300_splitterfromn300_4 , 0 , buf_n300_splitterfromn300_5 );
buf_AQFP buf_n308_n311_1_( clk_7 , n308 , 0 , buf_n308_n311_1 );
buf_AQFP buf_n308_n311_2_( clk_1 , buf_n308_n311_1 , 0 , buf_n308_n311_2 );
buf_AQFP buf_n309_n310_1_( clk_8 , n309 , 0 , buf_n309_n310_1 );
buf_AQFP buf_n311_splitterfromn311_1_( clk_5 , n311 , 0 , buf_n311_splitterfromn311_1 );
buf_AQFP buf_n311_splitterfromn311_2_( clk_7 , buf_n311_splitterfromn311_1 , 0 , buf_n311_splitterfromn311_2 );
buf_AQFP buf_n311_splitterfromn311_3_( clk_1 , buf_n311_splitterfromn311_2 , 0 , buf_n311_splitterfromn311_3 );
buf_AQFP buf_n312_splitterfromn312_1_( clk_7 , n312 , 0 , buf_n312_splitterfromn312_1 );
buf_AQFP buf_n312_splitterfromn312_2_( clk_1 , buf_n312_splitterfromn312_1 , 0 , buf_n312_splitterfromn312_2 );
buf_AQFP buf_n312_splitterfromn312_3_( clk_2 , buf_n312_splitterfromn312_2 , 0 , buf_n312_splitterfromn312_3 );
buf_AQFP buf_n312_splitterfromn312_4_( clk_3 , buf_n312_splitterfromn312_3 , 0 , buf_n312_splitterfromn312_4 );
buf_AQFP buf_splitterG1ton207n91_n207_1_( clk_7 , splitterG1ton207n91 , 0 , buf_splitterG1ton207n91_n207_1 );
buf_AQFP buf_splitterG1ton207n91_n207_2_( clk_1 , buf_splitterG1ton207n91_n207_1 , 0 , buf_splitterG1ton207n91_n207_2 );
buf_AQFP buf_splitterG1ton207n91_n207_3_( clk_3 , buf_splitterG1ton207n91_n207_2 , 0 , buf_splitterG1ton207n91_n207_3 );
buf_AQFP buf_splitterG1ton207n91_n207_4_( clk_5 , buf_splitterG1ton207n91_n207_3 , 0 , buf_splitterG1ton207n91_n207_4 );
buf_AQFP buf_splitterG1ton207n91_n207_5_( clk_7 , buf_splitterG1ton207n91_n207_4 , 0 , buf_splitterG1ton207n91_n207_5 );
buf_AQFP buf_splitterG1ton207n91_n207_6_( clk_1 , buf_splitterG1ton207n91_n207_5 , 0 , buf_splitterG1ton207n91_n207_6 );
buf_AQFP buf_splitterG1ton207n91_n207_7_( clk_3 , buf_splitterG1ton207n91_n207_6 , 0 , buf_splitterG1ton207n91_n207_7 );
buf_AQFP buf_splitterG1ton207n91_n207_8_( clk_5 , buf_splitterG1ton207n91_n207_7 , 0 , buf_splitterG1ton207n91_n207_8 );
buf_AQFP buf_splitterG1ton207n91_n207_9_( clk_7 , buf_splitterG1ton207n91_n207_8 , 0 , buf_splitterG1ton207n91_n207_9 );
buf_AQFP buf_splitterG1ton207n91_n207_10_( clk_1 , buf_splitterG1ton207n91_n207_9 , 0 , buf_splitterG1ton207n91_n207_10 );
buf_AQFP buf_splitterG1ton207n91_n207_11_( clk_2 , buf_splitterG1ton207n91_n207_10 , 0 , buf_splitterG1ton207n91_n207_11 );
buf_AQFP buf_splitterG1ton207n91_n207_12_( clk_4 , buf_splitterG1ton207n91_n207_11 , 0 , buf_splitterG1ton207n91_n207_12 );
buf_AQFP buf_splitterG1ton207n91_n208_1_( clk_7 , splitterG1ton207n91 , 0 , buf_splitterG1ton207n91_n208_1 );
buf_AQFP buf_splitterG1ton207n91_n208_2_( clk_1 , buf_splitterG1ton207n91_n208_1 , 0 , buf_splitterG1ton207n91_n208_2 );
buf_AQFP buf_splitterG1ton207n91_n208_3_( clk_3 , buf_splitterG1ton207n91_n208_2 , 0 , buf_splitterG1ton207n91_n208_3 );
buf_AQFP buf_splitterG1ton207n91_n208_4_( clk_5 , buf_splitterG1ton207n91_n208_3 , 0 , buf_splitterG1ton207n91_n208_4 );
buf_AQFP buf_splitterG1ton207n91_n208_5_( clk_7 , buf_splitterG1ton207n91_n208_4 , 0 , buf_splitterG1ton207n91_n208_5 );
buf_AQFP buf_splitterG1ton207n91_n208_6_( clk_1 , buf_splitterG1ton207n91_n208_5 , 0 , buf_splitterG1ton207n91_n208_6 );
buf_AQFP buf_splitterG1ton207n91_n208_7_( clk_3 , buf_splitterG1ton207n91_n208_6 , 0 , buf_splitterG1ton207n91_n208_7 );
buf_AQFP buf_splitterG1ton207n91_n208_8_( clk_5 , buf_splitterG1ton207n91_n208_7 , 0 , buf_splitterG1ton207n91_n208_8 );
buf_AQFP buf_splitterG1ton207n91_n208_9_( clk_7 , buf_splitterG1ton207n91_n208_8 , 0 , buf_splitterG1ton207n91_n208_9 );
buf_AQFP buf_splitterG1ton207n91_n208_10_( clk_1 , buf_splitterG1ton207n91_n208_9 , 0 , buf_splitterG1ton207n91_n208_10 );
buf_AQFP buf_splitterG1ton207n91_n208_11_( clk_3 , buf_splitterG1ton207n91_n208_10 , 0 , buf_splitterG1ton207n91_n208_11 );
buf_AQFP buf_splitterG1ton207n91_n208_12_( clk_5 , buf_splitterG1ton207n91_n208_11 , 0 , buf_splitterG1ton207n91_n208_12 );
buf_AQFP buf_splitterG10ton120n62_n120_1_( clk_4 , splitterG10ton120n62 , 0 , buf_splitterG10ton120n62_n120_1 );
buf_AQFP buf_splitterG10ton120n62_n121_1_( clk_4 , splitterG10ton120n62 , 0 , buf_splitterG10ton120n62_n121_1 );
buf_AQFP buf_splitterG10ton120n62_n223_1_( clk_4 , splitterG10ton120n62 , 0 , buf_splitterG10ton120n62_n223_1 );
buf_AQFP buf_splitterG10ton120n62_n223_2_( clk_6 , buf_splitterG10ton120n62_n223_1 , 0 , buf_splitterG10ton120n62_n223_2 );
buf_AQFP buf_splitterG10ton120n62_n223_3_( clk_8 , buf_splitterG10ton120n62_n223_2 , 0 , buf_splitterG10ton120n62_n223_3 );
buf_AQFP buf_splitterG10ton120n62_n223_4_( clk_2 , buf_splitterG10ton120n62_n223_3 , 0 , buf_splitterG10ton120n62_n223_4 );
buf_AQFP buf_splitterG10ton120n62_n223_5_( clk_4 , buf_splitterG10ton120n62_n223_4 , 0 , buf_splitterG10ton120n62_n223_5 );
buf_AQFP buf_splitterG10ton120n62_n223_6_( clk_6 , buf_splitterG10ton120n62_n223_5 , 0 , buf_splitterG10ton120n62_n223_6 );
buf_AQFP buf_splitterG10ton120n62_n223_7_( clk_8 , buf_splitterG10ton120n62_n223_6 , 0 , buf_splitterG10ton120n62_n223_7 );
buf_AQFP buf_splitterG10ton120n62_n223_8_( clk_2 , buf_splitterG10ton120n62_n223_7 , 0 , buf_splitterG10ton120n62_n223_8 );
buf_AQFP buf_splitterG10ton120n62_n223_9_( clk_4 , buf_splitterG10ton120n62_n223_8 , 0 , buf_splitterG10ton120n62_n223_9 );
buf_AQFP buf_splitterG10ton120n62_n223_10_( clk_6 , buf_splitterG10ton120n62_n223_9 , 0 , buf_splitterG10ton120n62_n223_10 );
buf_AQFP buf_splitterG10ton120n62_n223_11_( clk_8 , buf_splitterG10ton120n62_n223_10 , 0 , buf_splitterG10ton120n62_n223_11 );
buf_AQFP buf_splitterG10ton120n62_n223_12_( clk_2 , buf_splitterG10ton120n62_n223_11 , 0 , buf_splitterG10ton120n62_n223_12 );
buf_AQFP buf_splitterG10ton120n62_n223_13_( clk_4 , buf_splitterG10ton120n62_n223_12 , 0 , buf_splitterG10ton120n62_n223_13 );
buf_AQFP buf_splitterG10ton224n62_n224_1_( clk_5 , splitterG10ton224n62 , 0 , buf_splitterG10ton224n62_n224_1 );
buf_AQFP buf_splitterG10ton224n62_n224_2_( clk_7 , buf_splitterG10ton224n62_n224_1 , 0 , buf_splitterG10ton224n62_n224_2 );
buf_AQFP buf_splitterG10ton224n62_n224_3_( clk_1 , buf_splitterG10ton224n62_n224_2 , 0 , buf_splitterG10ton224n62_n224_3 );
buf_AQFP buf_splitterG10ton224n62_n224_4_( clk_3 , buf_splitterG10ton224n62_n224_3 , 0 , buf_splitterG10ton224n62_n224_4 );
buf_AQFP buf_splitterG10ton224n62_n224_5_( clk_5 , buf_splitterG10ton224n62_n224_4 , 0 , buf_splitterG10ton224n62_n224_5 );
buf_AQFP buf_splitterG10ton224n62_n224_6_( clk_7 , buf_splitterG10ton224n62_n224_5 , 0 , buf_splitterG10ton224n62_n224_6 );
buf_AQFP buf_splitterG10ton224n62_n224_7_( clk_1 , buf_splitterG10ton224n62_n224_6 , 0 , buf_splitterG10ton224n62_n224_7 );
buf_AQFP buf_splitterG10ton224n62_n224_8_( clk_3 , buf_splitterG10ton224n62_n224_7 , 0 , buf_splitterG10ton224n62_n224_8 );
buf_AQFP buf_splitterG10ton224n62_n224_9_( clk_5 , buf_splitterG10ton224n62_n224_8 , 0 , buf_splitterG10ton224n62_n224_9 );
buf_AQFP buf_splitterG10ton224n62_n224_10_( clk_7 , buf_splitterG10ton224n62_n224_9 , 0 , buf_splitterG10ton224n62_n224_10 );
buf_AQFP buf_splitterG10ton224n62_n224_11_( clk_1 , buf_splitterG10ton224n62_n224_10 , 0 , buf_splitterG10ton224n62_n224_11 );
buf_AQFP buf_splitterG10ton224n62_n224_12_( clk_2 , buf_splitterG10ton224n62_n224_11 , 0 , buf_splitterG10ton224n62_n224_12 );
buf_AQFP buf_splitterG10ton224n62_n224_13_( clk_4 , buf_splitterG10ton224n62_n224_12 , 0 , buf_splitterG10ton224n62_n224_13 );
buf_AQFP buf_splitterG11ton134n80_n255_1_( clk_4 , splitterG11ton134n80 , 0 , buf_splitterG11ton134n80_n255_1 );
buf_AQFP buf_splitterG11ton134n80_n255_2_( clk_6 , buf_splitterG11ton134n80_n255_1 , 0 , buf_splitterG11ton134n80_n255_2 );
buf_AQFP buf_splitterG11ton134n80_n255_3_( clk_8 , buf_splitterG11ton134n80_n255_2 , 0 , buf_splitterG11ton134n80_n255_3 );
buf_AQFP buf_splitterG11ton134n80_n255_4_( clk_2 , buf_splitterG11ton134n80_n255_3 , 0 , buf_splitterG11ton134n80_n255_4 );
buf_AQFP buf_splitterG11ton134n80_n255_5_( clk_4 , buf_splitterG11ton134n80_n255_4 , 0 , buf_splitterG11ton134n80_n255_5 );
buf_AQFP buf_splitterG11ton134n80_n255_6_( clk_6 , buf_splitterG11ton134n80_n255_5 , 0 , buf_splitterG11ton134n80_n255_6 );
buf_AQFP buf_splitterG11ton134n80_n255_7_( clk_8 , buf_splitterG11ton134n80_n255_6 , 0 , buf_splitterG11ton134n80_n255_7 );
buf_AQFP buf_splitterG11ton134n80_n255_8_( clk_2 , buf_splitterG11ton134n80_n255_7 , 0 , buf_splitterG11ton134n80_n255_8 );
buf_AQFP buf_splitterG11ton134n80_n255_9_( clk_4 , buf_splitterG11ton134n80_n255_8 , 0 , buf_splitterG11ton134n80_n255_9 );
buf_AQFP buf_splitterG11ton134n80_n255_10_( clk_6 , buf_splitterG11ton134n80_n255_9 , 0 , buf_splitterG11ton134n80_n255_10 );
buf_AQFP buf_splitterG11ton134n80_n255_11_( clk_8 , buf_splitterG11ton134n80_n255_10 , 0 , buf_splitterG11ton134n80_n255_11 );
buf_AQFP buf_splitterG11ton134n80_n255_12_( clk_2 , buf_splitterG11ton134n80_n255_11 , 0 , buf_splitterG11ton134n80_n255_12 );
buf_AQFP buf_splitterG11ton134n80_n255_13_( clk_4 , buf_splitterG11ton134n80_n255_12 , 0 , buf_splitterG11ton134n80_n255_13 );
buf_AQFP buf_splitterG11ton256n80_n256_1_( clk_5 , splitterG11ton256n80 , 0 , buf_splitterG11ton256n80_n256_1 );
buf_AQFP buf_splitterG11ton256n80_n256_2_( clk_7 , buf_splitterG11ton256n80_n256_1 , 0 , buf_splitterG11ton256n80_n256_2 );
buf_AQFP buf_splitterG11ton256n80_n256_3_( clk_1 , buf_splitterG11ton256n80_n256_2 , 0 , buf_splitterG11ton256n80_n256_3 );
buf_AQFP buf_splitterG11ton256n80_n256_4_( clk_3 , buf_splitterG11ton256n80_n256_3 , 0 , buf_splitterG11ton256n80_n256_4 );
buf_AQFP buf_splitterG11ton256n80_n256_5_( clk_5 , buf_splitterG11ton256n80_n256_4 , 0 , buf_splitterG11ton256n80_n256_5 );
buf_AQFP buf_splitterG11ton256n80_n256_6_( clk_7 , buf_splitterG11ton256n80_n256_5 , 0 , buf_splitterG11ton256n80_n256_6 );
buf_AQFP buf_splitterG11ton256n80_n256_7_( clk_1 , buf_splitterG11ton256n80_n256_6 , 0 , buf_splitterG11ton256n80_n256_7 );
buf_AQFP buf_splitterG11ton256n80_n256_8_( clk_3 , buf_splitterG11ton256n80_n256_7 , 0 , buf_splitterG11ton256n80_n256_8 );
buf_AQFP buf_splitterG11ton256n80_n256_9_( clk_5 , buf_splitterG11ton256n80_n256_8 , 0 , buf_splitterG11ton256n80_n256_9 );
buf_AQFP buf_splitterG11ton256n80_n256_10_( clk_7 , buf_splitterG11ton256n80_n256_9 , 0 , buf_splitterG11ton256n80_n256_10 );
buf_AQFP buf_splitterG11ton256n80_n256_11_( clk_1 , buf_splitterG11ton256n80_n256_10 , 0 , buf_splitterG11ton256n80_n256_11 );
buf_AQFP buf_splitterG11ton256n80_n256_12_( clk_3 , buf_splitterG11ton256n80_n256_11 , 0 , buf_splitterG11ton256n80_n256_12 );
buf_AQFP buf_splitterG11ton256n80_n256_13_( clk_4 , buf_splitterG11ton256n80_n256_12 , 0 , buf_splitterG11ton256n80_n256_13 );
buf_AQFP buf_splitterG12ton163n83_n258_1_( clk_7 , splitterG12ton163n83 , 0 , buf_splitterG12ton163n83_n258_1 );
buf_AQFP buf_splitterG12ton163n83_n258_2_( clk_1 , buf_splitterG12ton163n83_n258_1 , 0 , buf_splitterG12ton163n83_n258_2 );
buf_AQFP buf_splitterG12ton163n83_n258_3_( clk_3 , buf_splitterG12ton163n83_n258_2 , 0 , buf_splitterG12ton163n83_n258_3 );
buf_AQFP buf_splitterG12ton163n83_n258_4_( clk_5 , buf_splitterG12ton163n83_n258_3 , 0 , buf_splitterG12ton163n83_n258_4 );
buf_AQFP buf_splitterG12ton163n83_n258_5_( clk_7 , buf_splitterG12ton163n83_n258_4 , 0 , buf_splitterG12ton163n83_n258_5 );
buf_AQFP buf_splitterG12ton163n83_n258_6_( clk_1 , buf_splitterG12ton163n83_n258_5 , 0 , buf_splitterG12ton163n83_n258_6 );
buf_AQFP buf_splitterG12ton163n83_n258_7_( clk_3 , buf_splitterG12ton163n83_n258_6 , 0 , buf_splitterG12ton163n83_n258_7 );
buf_AQFP buf_splitterG12ton163n83_n258_8_( clk_5 , buf_splitterG12ton163n83_n258_7 , 0 , buf_splitterG12ton163n83_n258_8 );
buf_AQFP buf_splitterG12ton163n83_n258_9_( clk_7 , buf_splitterG12ton163n83_n258_8 , 0 , buf_splitterG12ton163n83_n258_9 );
buf_AQFP buf_splitterG12ton163n83_n258_10_( clk_1 , buf_splitterG12ton163n83_n258_9 , 0 , buf_splitterG12ton163n83_n258_10 );
buf_AQFP buf_splitterG12ton163n83_n258_11_( clk_3 , buf_splitterG12ton163n83_n258_10 , 0 , buf_splitterG12ton163n83_n258_11 );
buf_AQFP buf_splitterG12ton163n83_n258_12_( clk_4 , buf_splitterG12ton163n83_n258_11 , 0 , buf_splitterG12ton163n83_n258_12 );
buf_AQFP buf_splitterG12ton163n83_n258_13_( clk_5 , buf_splitterG12ton163n83_n258_12 , 0 , buf_splitterG12ton163n83_n258_13 );
buf_AQFP buf_splitterG12ton259n83_n259_1_( clk_8 , splitterG12ton259n83 , 0 , buf_splitterG12ton259n83_n259_1 );
buf_AQFP buf_splitterG12ton259n83_n259_2_( clk_2 , buf_splitterG12ton259n83_n259_1 , 0 , buf_splitterG12ton259n83_n259_2 );
buf_AQFP buf_splitterG12ton259n83_n259_3_( clk_4 , buf_splitterG12ton259n83_n259_2 , 0 , buf_splitterG12ton259n83_n259_3 );
buf_AQFP buf_splitterG12ton259n83_n259_4_( clk_6 , buf_splitterG12ton259n83_n259_3 , 0 , buf_splitterG12ton259n83_n259_4 );
buf_AQFP buf_splitterG12ton259n83_n259_5_( clk_8 , buf_splitterG12ton259n83_n259_4 , 0 , buf_splitterG12ton259n83_n259_5 );
buf_AQFP buf_splitterG12ton259n83_n259_6_( clk_2 , buf_splitterG12ton259n83_n259_5 , 0 , buf_splitterG12ton259n83_n259_6 );
buf_AQFP buf_splitterG12ton259n83_n259_7_( clk_4 , buf_splitterG12ton259n83_n259_6 , 0 , buf_splitterG12ton259n83_n259_7 );
buf_AQFP buf_splitterG12ton259n83_n259_8_( clk_6 , buf_splitterG12ton259n83_n259_7 , 0 , buf_splitterG12ton259n83_n259_8 );
buf_AQFP buf_splitterG12ton259n83_n259_9_( clk_8 , buf_splitterG12ton259n83_n259_8 , 0 , buf_splitterG12ton259n83_n259_9 );
buf_AQFP buf_splitterG12ton259n83_n259_10_( clk_1 , buf_splitterG12ton259n83_n259_9 , 0 , buf_splitterG12ton259n83_n259_10 );
buf_AQFP buf_splitterG12ton259n83_n259_11_( clk_3 , buf_splitterG12ton259n83_n259_10 , 0 , buf_splitterG12ton259n83_n259_11 );
buf_AQFP buf_splitterG12ton259n83_n259_12_( clk_5 , buf_splitterG12ton259n83_n259_11 , 0 , buf_splitterG12ton259n83_n259_12 );
buf_AQFP buf_splitterG13ton111n80_n111_1_( clk_4 , splitterG13ton111n80 , 0 , buf_splitterG13ton111n80_n111_1 );
buf_AQFP buf_splitterG13ton111n80_n111_2_( clk_6 , buf_splitterG13ton111n80_n111_1 , 0 , buf_splitterG13ton111n80_n111_2 );
buf_AQFP buf_splitterG13ton111n80_n112_1_( clk_4 , splitterG13ton111n80 , 0 , buf_splitterG13ton111n80_n112_1 );
buf_AQFP buf_splitterG13ton111n80_n112_2_( clk_6 , buf_splitterG13ton111n80_n112_1 , 0 , buf_splitterG13ton111n80_n112_2 );
buf_AQFP buf_splitterG13ton111n80_n261_1_( clk_4 , splitterG13ton111n80 , 0 , buf_splitterG13ton111n80_n261_1 );
buf_AQFP buf_splitterG13ton111n80_n261_2_( clk_6 , buf_splitterG13ton111n80_n261_1 , 0 , buf_splitterG13ton111n80_n261_2 );
buf_AQFP buf_splitterG13ton111n80_n261_3_( clk_8 , buf_splitterG13ton111n80_n261_2 , 0 , buf_splitterG13ton111n80_n261_3 );
buf_AQFP buf_splitterG13ton111n80_n261_4_( clk_2 , buf_splitterG13ton111n80_n261_3 , 0 , buf_splitterG13ton111n80_n261_4 );
buf_AQFP buf_splitterG13ton111n80_n261_5_( clk_4 , buf_splitterG13ton111n80_n261_4 , 0 , buf_splitterG13ton111n80_n261_5 );
buf_AQFP buf_splitterG13ton111n80_n261_6_( clk_6 , buf_splitterG13ton111n80_n261_5 , 0 , buf_splitterG13ton111n80_n261_6 );
buf_AQFP buf_splitterG13ton111n80_n261_7_( clk_8 , buf_splitterG13ton111n80_n261_6 , 0 , buf_splitterG13ton111n80_n261_7 );
buf_AQFP buf_splitterG13ton111n80_n261_8_( clk_2 , buf_splitterG13ton111n80_n261_7 , 0 , buf_splitterG13ton111n80_n261_8 );
buf_AQFP buf_splitterG13ton111n80_n261_9_( clk_3 , buf_splitterG13ton111n80_n261_8 , 0 , buf_splitterG13ton111n80_n261_9 );
buf_AQFP buf_splitterG13ton111n80_n261_10_( clk_5 , buf_splitterG13ton111n80_n261_9 , 0 , buf_splitterG13ton111n80_n261_10 );
buf_AQFP buf_splitterG13ton111n80_n261_11_( clk_7 , buf_splitterG13ton111n80_n261_10 , 0 , buf_splitterG13ton111n80_n261_11 );
buf_AQFP buf_splitterG13ton111n80_n261_12_( clk_1 , buf_splitterG13ton111n80_n261_11 , 0 , buf_splitterG13ton111n80_n261_12 );
buf_AQFP buf_splitterG13ton111n80_n261_13_( clk_3 , buf_splitterG13ton111n80_n261_12 , 0 , buf_splitterG13ton111n80_n261_13 );
buf_AQFP buf_splitterG13ton111n80_n261_14_( clk_5 , buf_splitterG13ton111n80_n261_13 , 0 , buf_splitterG13ton111n80_n261_14 );
buf_AQFP buf_splitterG13ton111n80_n261_15_( clk_7 , buf_splitterG13ton111n80_n261_14 , 0 , buf_splitterG13ton111n80_n261_15 );
buf_AQFP buf_splitterG13ton262n80_n262_1_( clk_5 , splitterG13ton262n80 , 0 , buf_splitterG13ton262n80_n262_1 );
buf_AQFP buf_splitterG13ton262n80_n262_2_( clk_7 , buf_splitterG13ton262n80_n262_1 , 0 , buf_splitterG13ton262n80_n262_2 );
buf_AQFP buf_splitterG13ton262n80_n262_3_( clk_1 , buf_splitterG13ton262n80_n262_2 , 0 , buf_splitterG13ton262n80_n262_3 );
buf_AQFP buf_splitterG13ton262n80_n262_4_( clk_3 , buf_splitterG13ton262n80_n262_3 , 0 , buf_splitterG13ton262n80_n262_4 );
buf_AQFP buf_splitterG13ton262n80_n262_5_( clk_5 , buf_splitterG13ton262n80_n262_4 , 0 , buf_splitterG13ton262n80_n262_5 );
buf_AQFP buf_splitterG13ton262n80_n262_6_( clk_7 , buf_splitterG13ton262n80_n262_5 , 0 , buf_splitterG13ton262n80_n262_6 );
buf_AQFP buf_splitterG13ton262n80_n262_7_( clk_1 , buf_splitterG13ton262n80_n262_6 , 0 , buf_splitterG13ton262n80_n262_7 );
buf_AQFP buf_splitterG13ton262n80_n262_8_( clk_3 , buf_splitterG13ton262n80_n262_7 , 0 , buf_splitterG13ton262n80_n262_8 );
buf_AQFP buf_splitterG13ton262n80_n262_9_( clk_5 , buf_splitterG13ton262n80_n262_8 , 0 , buf_splitterG13ton262n80_n262_9 );
buf_AQFP buf_splitterG13ton262n80_n262_10_( clk_7 , buf_splitterG13ton262n80_n262_9 , 0 , buf_splitterG13ton262n80_n262_10 );
buf_AQFP buf_splitterG13ton262n80_n262_11_( clk_1 , buf_splitterG13ton262n80_n262_10 , 0 , buf_splitterG13ton262n80_n262_11 );
buf_AQFP buf_splitterG13ton262n80_n262_12_( clk_3 , buf_splitterG13ton262n80_n262_11 , 0 , buf_splitterG13ton262n80_n262_12 );
buf_AQFP buf_splitterG13ton262n80_n262_13_( clk_5 , buf_splitterG13ton262n80_n262_12 , 0 , buf_splitterG13ton262n80_n262_13 );
buf_AQFP buf_splitterG13ton262n80_n262_14_( clk_6 , buf_splitterG13ton262n80_n262_13 , 0 , buf_splitterG13ton262n80_n262_14 );
buf_AQFP buf_splitterG14ton103n265_n180_1_( clk_3 , splitterG14ton103n265 , 0 , buf_splitterG14ton103n265_n180_1 );
buf_AQFP buf_splitterG14ton181n265_n264_1_( clk_7 , splitterG14ton181n265 , 0 , buf_splitterG14ton181n265_n264_1 );
buf_AQFP buf_splitterG14ton181n265_n264_2_( clk_1 , buf_splitterG14ton181n265_n264_1 , 0 , buf_splitterG14ton181n265_n264_2 );
buf_AQFP buf_splitterG14ton181n265_n264_3_( clk_3 , buf_splitterG14ton181n265_n264_2 , 0 , buf_splitterG14ton181n265_n264_3 );
buf_AQFP buf_splitterG14ton181n265_n264_4_( clk_5 , buf_splitterG14ton181n265_n264_3 , 0 , buf_splitterG14ton181n265_n264_4 );
buf_AQFP buf_splitterG14ton181n265_n264_5_( clk_6 , buf_splitterG14ton181n265_n264_4 , 0 , buf_splitterG14ton181n265_n264_5 );
buf_AQFP buf_splitterG14ton181n265_n264_6_( clk_7 , buf_splitterG14ton181n265_n264_5 , 0 , buf_splitterG14ton181n265_n264_6 );
buf_AQFP buf_splitterG14ton181n265_n264_7_( clk_1 , buf_splitterG14ton181n265_n264_6 , 0 , buf_splitterG14ton181n265_n264_7 );
buf_AQFP buf_splitterG14ton181n265_n264_8_( clk_3 , buf_splitterG14ton181n265_n264_7 , 0 , buf_splitterG14ton181n265_n264_8 );
buf_AQFP buf_splitterG14ton181n265_n264_9_( clk_5 , buf_splitterG14ton181n265_n264_8 , 0 , buf_splitterG14ton181n265_n264_9 );
buf_AQFP buf_splitterG14ton181n265_n264_10_( clk_7 , buf_splitterG14ton181n265_n264_9 , 0 , buf_splitterG14ton181n265_n264_10 );
buf_AQFP buf_splitterG14ton181n265_n264_11_( clk_1 , buf_splitterG14ton181n265_n264_10 , 0 , buf_splitterG14ton181n265_n264_11 );
buf_AQFP buf_splitterG14ton181n265_n264_12_( clk_3 , buf_splitterG14ton181n265_n264_11 , 0 , buf_splitterG14ton181n265_n264_12 );
buf_AQFP buf_splitterG14ton181n265_n264_13_( clk_5 , buf_splitterG14ton181n265_n264_12 , 0 , buf_splitterG14ton181n265_n264_13 );
buf_AQFP buf_splitterG14ton181n265_n265_1_( clk_7 , splitterG14ton181n265 , 0 , buf_splitterG14ton181n265_n265_1 );
buf_AQFP buf_splitterG14ton181n265_n265_2_( clk_1 , buf_splitterG14ton181n265_n265_1 , 0 , buf_splitterG14ton181n265_n265_2 );
buf_AQFP buf_splitterG14ton181n265_n265_3_( clk_3 , buf_splitterG14ton181n265_n265_2 , 0 , buf_splitterG14ton181n265_n265_3 );
buf_AQFP buf_splitterG14ton181n265_n265_4_( clk_5 , buf_splitterG14ton181n265_n265_3 , 0 , buf_splitterG14ton181n265_n265_4 );
buf_AQFP buf_splitterG14ton181n265_n265_5_( clk_7 , buf_splitterG14ton181n265_n265_4 , 0 , buf_splitterG14ton181n265_n265_5 );
buf_AQFP buf_splitterG14ton181n265_n265_6_( clk_1 , buf_splitterG14ton181n265_n265_5 , 0 , buf_splitterG14ton181n265_n265_6 );
buf_AQFP buf_splitterG14ton181n265_n265_7_( clk_3 , buf_splitterG14ton181n265_n265_6 , 0 , buf_splitterG14ton181n265_n265_7 );
buf_AQFP buf_splitterG14ton181n265_n265_8_( clk_5 , buf_splitterG14ton181n265_n265_7 , 0 , buf_splitterG14ton181n265_n265_8 );
buf_AQFP buf_splitterG14ton181n265_n265_9_( clk_7 , buf_splitterG14ton181n265_n265_8 , 0 , buf_splitterG14ton181n265_n265_9 );
buf_AQFP buf_splitterG14ton181n265_n265_10_( clk_1 , buf_splitterG14ton181n265_n265_9 , 0 , buf_splitterG14ton181n265_n265_10 );
buf_AQFP buf_splitterG14ton181n265_n265_11_( clk_2 , buf_splitterG14ton181n265_n265_10 , 0 , buf_splitterG14ton181n265_n265_11 );
buf_AQFP buf_splitterG14ton181n265_n265_12_( clk_4 , buf_splitterG14ton181n265_n265_11 , 0 , buf_splitterG14ton181n265_n265_12 );
buf_AQFP buf_splitterG14ton181n265_n265_13_( clk_5 , buf_splitterG14ton181n265_n265_12 , 0 , buf_splitterG14ton181n265_n265_13 );
buf_AQFP buf_splitterG15ton134n62_n226_1_( clk_4 , splitterG15ton134n62 , 0 , buf_splitterG15ton134n62_n226_1 );
buf_AQFP buf_splitterG15ton134n62_n226_2_( clk_6 , buf_splitterG15ton134n62_n226_1 , 0 , buf_splitterG15ton134n62_n226_2 );
buf_AQFP buf_splitterG15ton134n62_n226_3_( clk_8 , buf_splitterG15ton134n62_n226_2 , 0 , buf_splitterG15ton134n62_n226_3 );
buf_AQFP buf_splitterG15ton134n62_n226_4_( clk_2 , buf_splitterG15ton134n62_n226_3 , 0 , buf_splitterG15ton134n62_n226_4 );
buf_AQFP buf_splitterG15ton134n62_n226_5_( clk_4 , buf_splitterG15ton134n62_n226_4 , 0 , buf_splitterG15ton134n62_n226_5 );
buf_AQFP buf_splitterG15ton134n62_n226_6_( clk_6 , buf_splitterG15ton134n62_n226_5 , 0 , buf_splitterG15ton134n62_n226_6 );
buf_AQFP buf_splitterG15ton134n62_n226_7_( clk_8 , buf_splitterG15ton134n62_n226_6 , 0 , buf_splitterG15ton134n62_n226_7 );
buf_AQFP buf_splitterG15ton134n62_n226_8_( clk_2 , buf_splitterG15ton134n62_n226_7 , 0 , buf_splitterG15ton134n62_n226_8 );
buf_AQFP buf_splitterG15ton134n62_n226_9_( clk_4 , buf_splitterG15ton134n62_n226_8 , 0 , buf_splitterG15ton134n62_n226_9 );
buf_AQFP buf_splitterG15ton134n62_n226_10_( clk_6 , buf_splitterG15ton134n62_n226_9 , 0 , buf_splitterG15ton134n62_n226_10 );
buf_AQFP buf_splitterG15ton134n62_n226_11_( clk_8 , buf_splitterG15ton134n62_n226_10 , 0 , buf_splitterG15ton134n62_n226_11 );
buf_AQFP buf_splitterG15ton134n62_n226_12_( clk_1 , buf_splitterG15ton134n62_n226_11 , 0 , buf_splitterG15ton134n62_n226_12 );
buf_AQFP buf_splitterG15ton134n62_n226_13_( clk_3 , buf_splitterG15ton134n62_n226_12 , 0 , buf_splitterG15ton134n62_n226_13 );
buf_AQFP buf_splitterG15ton134n62_n226_14_( clk_5 , buf_splitterG15ton134n62_n226_13 , 0 , buf_splitterG15ton134n62_n226_14 );
buf_AQFP buf_splitterG15ton227n62_n227_1_( clk_5 , splitterG15ton227n62 , 0 , buf_splitterG15ton227n62_n227_1 );
buf_AQFP buf_splitterG15ton227n62_n227_2_( clk_7 , buf_splitterG15ton227n62_n227_1 , 0 , buf_splitterG15ton227n62_n227_2 );
buf_AQFP buf_splitterG15ton227n62_n227_3_( clk_1 , buf_splitterG15ton227n62_n227_2 , 0 , buf_splitterG15ton227n62_n227_3 );
buf_AQFP buf_splitterG15ton227n62_n227_4_( clk_3 , buf_splitterG15ton227n62_n227_3 , 0 , buf_splitterG15ton227n62_n227_4 );
buf_AQFP buf_splitterG15ton227n62_n227_5_( clk_5 , buf_splitterG15ton227n62_n227_4 , 0 , buf_splitterG15ton227n62_n227_5 );
buf_AQFP buf_splitterG15ton227n62_n227_6_( clk_7 , buf_splitterG15ton227n62_n227_5 , 0 , buf_splitterG15ton227n62_n227_6 );
buf_AQFP buf_splitterG15ton227n62_n227_7_( clk_1 , buf_splitterG15ton227n62_n227_6 , 0 , buf_splitterG15ton227n62_n227_7 );
buf_AQFP buf_splitterG15ton227n62_n227_8_( clk_3 , buf_splitterG15ton227n62_n227_7 , 0 , buf_splitterG15ton227n62_n227_8 );
buf_AQFP buf_splitterG15ton227n62_n227_9_( clk_5 , buf_splitterG15ton227n62_n227_8 , 0 , buf_splitterG15ton227n62_n227_9 );
buf_AQFP buf_splitterG15ton227n62_n227_10_( clk_7 , buf_splitterG15ton227n62_n227_9 , 0 , buf_splitterG15ton227n62_n227_10 );
buf_AQFP buf_splitterG15ton227n62_n227_11_( clk_1 , buf_splitterG15ton227n62_n227_10 , 0 , buf_splitterG15ton227n62_n227_11 );
buf_AQFP buf_splitterG15ton227n62_n227_12_( clk_3 , buf_splitterG15ton227n62_n227_11 , 0 , buf_splitterG15ton227n62_n227_12 );
buf_AQFP buf_splitterG15ton227n62_n227_13_( clk_5 , buf_splitterG15ton227n62_n227_12 , 0 , buf_splitterG15ton227n62_n227_13 );
buf_AQFP buf_splitterG15ton227n62_n227_14_( clk_7 , buf_splitterG15ton227n62_n227_13 , 0 , buf_splitterG15ton227n62_n227_14 );
buf_AQFP buf_splitterG16ton106n65_n229_1_( clk_7 , splitterG16ton106n65 , 0 , buf_splitterG16ton106n65_n229_1 );
buf_AQFP buf_splitterG16ton106n65_n229_2_( clk_1 , buf_splitterG16ton106n65_n229_1 , 0 , buf_splitterG16ton106n65_n229_2 );
buf_AQFP buf_splitterG16ton106n65_n229_3_( clk_3 , buf_splitterG16ton106n65_n229_2 , 0 , buf_splitterG16ton106n65_n229_3 );
buf_AQFP buf_splitterG16ton106n65_n229_4_( clk_5 , buf_splitterG16ton106n65_n229_3 , 0 , buf_splitterG16ton106n65_n229_4 );
buf_AQFP buf_splitterG16ton106n65_n229_5_( clk_7 , buf_splitterG16ton106n65_n229_4 , 0 , buf_splitterG16ton106n65_n229_5 );
buf_AQFP buf_splitterG16ton106n65_n229_6_( clk_1 , buf_splitterG16ton106n65_n229_5 , 0 , buf_splitterG16ton106n65_n229_6 );
buf_AQFP buf_splitterG16ton106n65_n229_7_( clk_2 , buf_splitterG16ton106n65_n229_6 , 0 , buf_splitterG16ton106n65_n229_7 );
buf_AQFP buf_splitterG16ton106n65_n229_8_( clk_4 , buf_splitterG16ton106n65_n229_7 , 0 , buf_splitterG16ton106n65_n229_8 );
buf_AQFP buf_splitterG16ton106n65_n229_9_( clk_6 , buf_splitterG16ton106n65_n229_8 , 0 , buf_splitterG16ton106n65_n229_9 );
buf_AQFP buf_splitterG16ton106n65_n229_10_( clk_8 , buf_splitterG16ton106n65_n229_9 , 0 , buf_splitterG16ton106n65_n229_10 );
buf_AQFP buf_splitterG16ton106n65_n229_11_( clk_2 , buf_splitterG16ton106n65_n229_10 , 0 , buf_splitterG16ton106n65_n229_11 );
buf_AQFP buf_splitterG16ton106n65_n229_12_( clk_4 , buf_splitterG16ton106n65_n229_11 , 0 , buf_splitterG16ton106n65_n229_12 );
buf_AQFP buf_splitterG16ton106n65_n229_13_( clk_6 , buf_splitterG16ton106n65_n229_12 , 0 , buf_splitterG16ton106n65_n229_13 );
buf_AQFP buf_splitterG16ton230n65_n230_1_( clk_8 , splitterG16ton230n65 , 0 , buf_splitterG16ton230n65_n230_1 );
buf_AQFP buf_splitterG16ton230n65_n230_2_( clk_2 , buf_splitterG16ton230n65_n230_1 , 0 , buf_splitterG16ton230n65_n230_2 );
buf_AQFP buf_splitterG16ton230n65_n230_3_( clk_4 , buf_splitterG16ton230n65_n230_2 , 0 , buf_splitterG16ton230n65_n230_3 );
buf_AQFP buf_splitterG16ton230n65_n230_4_( clk_6 , buf_splitterG16ton230n65_n230_3 , 0 , buf_splitterG16ton230n65_n230_4 );
buf_AQFP buf_splitterG16ton230n65_n230_5_( clk_8 , buf_splitterG16ton230n65_n230_4 , 0 , buf_splitterG16ton230n65_n230_5 );
buf_AQFP buf_splitterG16ton230n65_n230_6_( clk_2 , buf_splitterG16ton230n65_n230_5 , 0 , buf_splitterG16ton230n65_n230_6 );
buf_AQFP buf_splitterG16ton230n65_n230_7_( clk_4 , buf_splitterG16ton230n65_n230_6 , 0 , buf_splitterG16ton230n65_n230_7 );
buf_AQFP buf_splitterG16ton230n65_n230_8_( clk_6 , buf_splitterG16ton230n65_n230_7 , 0 , buf_splitterG16ton230n65_n230_8 );
buf_AQFP buf_splitterG16ton230n65_n230_9_( clk_8 , buf_splitterG16ton230n65_n230_8 , 0 , buf_splitterG16ton230n65_n230_9 );
buf_AQFP buf_splitterG16ton230n65_n230_10_( clk_2 , buf_splitterG16ton230n65_n230_9 , 0 , buf_splitterG16ton230n65_n230_10 );
buf_AQFP buf_splitterG16ton230n65_n230_11_( clk_4 , buf_splitterG16ton230n65_n230_10 , 0 , buf_splitterG16ton230n65_n230_11 );
buf_AQFP buf_splitterG16ton230n65_n230_12_( clk_6 , buf_splitterG16ton230n65_n230_11 , 0 , buf_splitterG16ton230n65_n230_12 );
buf_AQFP buf_splitterfromG17_n74_1_( clk_6 , splitterfromG17 , 0 , buf_splitterfromG17_n74_1 );
buf_AQFP buf_splitterfromG17_n74_2_( clk_8 , buf_splitterfromG17_n74_1 , 0 , buf_splitterfromG17_n74_2 );
buf_AQFP buf_splitterfromG17_n74_3_( clk_2 , buf_splitterfromG17_n74_2 , 0 , buf_splitterfromG17_n74_3 );
buf_AQFP buf_splitterfromG17_n74_4_( clk_4 , buf_splitterfromG17_n74_3 , 0 , buf_splitterfromG17_n74_4 );
buf_AQFP buf_splitterfromG17_n74_5_( clk_5 , buf_splitterfromG17_n74_4 , 0 , buf_splitterfromG17_n74_5 );
buf_AQFP buf_splitterfromG18_n35_1_( clk_7 , splitterfromG18 , 0 , buf_splitterfromG18_n35_1 );
buf_AQFP buf_splitterfromG18_n35_2_( clk_1 , buf_splitterfromG18_n35_1 , 0 , buf_splitterfromG18_n35_2 );
buf_AQFP buf_splitterfromG18_n35_3_( clk_3 , buf_splitterfromG18_n35_2 , 0 , buf_splitterfromG18_n35_3 );
buf_AQFP buf_splitterfromG19_n128_1_( clk_8 , splitterfromG19 , 0 , buf_splitterfromG19_n128_1 );
buf_AQFP buf_splitterfromG19_n128_2_( clk_2 , buf_splitterfromG19_n128_1 , 0 , buf_splitterfromG19_n128_2 );
buf_AQFP buf_splitterfromG19_n128_3_( clk_4 , buf_splitterfromG19_n128_2 , 0 , buf_splitterfromG19_n128_3 );
buf_AQFP buf_splitterfromG19_n128_4_( clk_6 , buf_splitterfromG19_n128_3 , 0 , buf_splitterfromG19_n128_4 );
buf_AQFP buf_splitterfromG19_n128_5_( clk_7 , buf_splitterfromG19_n128_4 , 0 , buf_splitterfromG19_n128_5 );
buf_AQFP buf_splitterG2ton146n46_n146_1_( clk_4 , splitterG2ton146n46 , 0 , buf_splitterG2ton146n46_n146_1 );
buf_AQFP buf_splitterG2ton146n46_n147_1_( clk_4 , splitterG2ton146n46 , 0 , buf_splitterG2ton146n46_n147_1 );
buf_AQFP buf_splitterG2ton146n46_n210_1_( clk_4 , splitterG2ton146n46 , 0 , buf_splitterG2ton146n46_n210_1 );
buf_AQFP buf_splitterG2ton146n46_n210_2_( clk_6 , buf_splitterG2ton146n46_n210_1 , 0 , buf_splitterG2ton146n46_n210_2 );
buf_AQFP buf_splitterG2ton146n46_n210_3_( clk_8 , buf_splitterG2ton146n46_n210_2 , 0 , buf_splitterG2ton146n46_n210_3 );
buf_AQFP buf_splitterG2ton146n46_n210_4_( clk_2 , buf_splitterG2ton146n46_n210_3 , 0 , buf_splitterG2ton146n46_n210_4 );
buf_AQFP buf_splitterG2ton146n46_n210_5_( clk_4 , buf_splitterG2ton146n46_n210_4 , 0 , buf_splitterG2ton146n46_n210_5 );
buf_AQFP buf_splitterG2ton146n46_n210_6_( clk_6 , buf_splitterG2ton146n46_n210_5 , 0 , buf_splitterG2ton146n46_n210_6 );
buf_AQFP buf_splitterG2ton146n46_n210_7_( clk_8 , buf_splitterG2ton146n46_n210_6 , 0 , buf_splitterG2ton146n46_n210_7 );
buf_AQFP buf_splitterG2ton146n46_n210_8_( clk_2 , buf_splitterG2ton146n46_n210_7 , 0 , buf_splitterG2ton146n46_n210_8 );
buf_AQFP buf_splitterG2ton146n46_n210_9_( clk_4 , buf_splitterG2ton146n46_n210_8 , 0 , buf_splitterG2ton146n46_n210_9 );
buf_AQFP buf_splitterG2ton146n46_n210_10_( clk_6 , buf_splitterG2ton146n46_n210_9 , 0 , buf_splitterG2ton146n46_n210_10 );
buf_AQFP buf_splitterG2ton146n46_n210_11_( clk_8 , buf_splitterG2ton146n46_n210_10 , 0 , buf_splitterG2ton146n46_n210_11 );
buf_AQFP buf_splitterG2ton146n46_n210_12_( clk_2 , buf_splitterG2ton146n46_n210_11 , 0 , buf_splitterG2ton146n46_n210_12 );
buf_AQFP buf_splitterG2ton146n46_n210_13_( clk_4 , buf_splitterG2ton146n46_n210_12 , 0 , buf_splitterG2ton146n46_n210_13 );
buf_AQFP buf_splitterG2ton146n46_n210_14_( clk_6 , buf_splitterG2ton146n46_n210_13 , 0 , buf_splitterG2ton146n46_n210_14 );
buf_AQFP buf_splitterG2ton211n46_n211_1_( clk_5 , splitterG2ton211n46 , 0 , buf_splitterG2ton211n46_n211_1 );
buf_AQFP buf_splitterG2ton211n46_n211_2_( clk_7 , buf_splitterG2ton211n46_n211_1 , 0 , buf_splitterG2ton211n46_n211_2 );
buf_AQFP buf_splitterG2ton211n46_n211_3_( clk_1 , buf_splitterG2ton211n46_n211_2 , 0 , buf_splitterG2ton211n46_n211_3 );
buf_AQFP buf_splitterG2ton211n46_n211_4_( clk_3 , buf_splitterG2ton211n46_n211_3 , 0 , buf_splitterG2ton211n46_n211_4 );
buf_AQFP buf_splitterG2ton211n46_n211_5_( clk_5 , buf_splitterG2ton211n46_n211_4 , 0 , buf_splitterG2ton211n46_n211_5 );
buf_AQFP buf_splitterG2ton211n46_n211_6_( clk_7 , buf_splitterG2ton211n46_n211_5 , 0 , buf_splitterG2ton211n46_n211_6 );
buf_AQFP buf_splitterG2ton211n46_n211_7_( clk_1 , buf_splitterG2ton211n46_n211_6 , 0 , buf_splitterG2ton211n46_n211_7 );
buf_AQFP buf_splitterG2ton211n46_n211_8_( clk_3 , buf_splitterG2ton211n46_n211_7 , 0 , buf_splitterG2ton211n46_n211_8 );
buf_AQFP buf_splitterG2ton211n46_n211_9_( clk_5 , buf_splitterG2ton211n46_n211_8 , 0 , buf_splitterG2ton211n46_n211_9 );
buf_AQFP buf_splitterG2ton211n46_n211_10_( clk_7 , buf_splitterG2ton211n46_n211_9 , 0 , buf_splitterG2ton211n46_n211_10 );
buf_AQFP buf_splitterG2ton211n46_n211_11_( clk_1 , buf_splitterG2ton211n46_n211_10 , 0 , buf_splitterG2ton211n46_n211_11 );
buf_AQFP buf_splitterG2ton211n46_n211_12_( clk_3 , buf_splitterG2ton211n46_n211_11 , 0 , buf_splitterG2ton211n46_n211_12 );
buf_AQFP buf_splitterG2ton211n46_n211_13_( clk_5 , buf_splitterG2ton211n46_n211_12 , 0 , buf_splitterG2ton211n46_n211_13 );
buf_AQFP buf_splitterG2ton211n46_n211_14_( clk_7 , buf_splitterG2ton211n46_n211_13 , 0 , buf_splitterG2ton211n46_n211_14 );
buf_AQFP buf_splitterfromG20_n178_1_( clk_6 , splitterfromG20 , 0 , buf_splitterfromG20_n178_1 );
buf_AQFP buf_splitterfromG20_n178_2_( clk_7 , buf_splitterfromG20_n178_1 , 0 , buf_splitterfromG20_n178_2 );
buf_AQFP buf_splitterfromG20_n178_3_( clk_1 , buf_splitterfromG20_n178_2 , 0 , buf_splitterfromG20_n178_3 );
buf_AQFP buf_splitterfromG20_n178_4_( clk_3 , buf_splitterfromG20_n178_3 , 0 , buf_splitterfromG20_n178_4 );
buf_AQFP buf_splitterfromG20_n178_5_( clk_4 , buf_splitterfromG20_n178_4 , 0 , buf_splitterfromG20_n178_5 );
buf_AQFP buf_splitterfromG20_n178_6_( clk_6 , buf_splitterfromG20_n178_5 , 0 , buf_splitterfromG20_n178_6 );
buf_AQFP buf_splitterG23ton109n200_n127_1_( clk_5 , splitterG23ton109n200 , 0 , buf_splitterG23ton109n200_n127_1 );
buf_AQFP buf_splitterG23ton109n200_n127_2_( clk_7 , buf_splitterG23ton109n200_n127_1 , 0 , buf_splitterG23ton109n200_n127_2 );
buf_AQFP buf_splitterG23ton109n200_n127_3_( clk_1 , buf_splitterG23ton109n200_n127_2 , 0 , buf_splitterG23ton109n200_n127_3 );
buf_AQFP buf_splitterG23ton109n200_n127_4_( clk_3 , buf_splitterG23ton109n200_n127_3 , 0 , buf_splitterG23ton109n200_n127_4 );
buf_AQFP buf_splitterG23ton109n200_n200_1_( clk_4 , splitterG23ton109n200 , 0 , buf_splitterG23ton109n200_n200_1 );
buf_AQFP buf_splitterG24ton200n88_n200_1_( clk_5 , splitterG24ton200n88 , 0 , buf_splitterG24ton200n88_n200_1 );
buf_AQFP buf_splitterG24ton200n88_n34_1_( clk_4 , splitterG24ton200n88 , 0 , buf_splitterG24ton200n88_n34_1 );
buf_AQFP buf_splitterG24ton200n88_n34_2_( clk_5 , buf_splitterG24ton200n88_n34_1 , 0 , buf_splitterG24ton200n88_n34_2 );
buf_AQFP buf_splitterG24ton200n88_n34_3_( clk_6 , buf_splitterG24ton200n88_n34_2 , 0 , buf_splitterG24ton200n88_n34_3 );
buf_AQFP buf_splitterG24ton200n88_n34_4_( clk_8 , buf_splitterG24ton200n88_n34_3 , 0 , buf_splitterG24ton200n88_n34_4 );
buf_AQFP buf_splitterG24ton200n88_n34_5_( clk_2 , buf_splitterG24ton200n88_n34_4 , 0 , buf_splitterG24ton200n88_n34_5 );
buf_AQFP buf_splitterG25ton193n281_n281_1_( clk_4 , splitterG25ton193n281 , 0 , buf_splitterG25ton193n281_n281_1 );
buf_AQFP buf_splitterG25ton193n281_n281_2_( clk_5 , buf_splitterG25ton193n281_n281_1 , 0 , buf_splitterG25ton193n281_n281_2 );
buf_AQFP buf_splitterG25ton193n281_n281_3_( clk_6 , buf_splitterG25ton193n281_n281_2 , 0 , buf_splitterG25ton193n281_n281_3 );
buf_AQFP buf_splitterG25ton193n281_n281_4_( clk_8 , buf_splitterG25ton193n281_n281_3 , 0 , buf_splitterG25ton193n281_n281_4 );
buf_AQFP buf_splitterG25ton193n281_n281_5_( clk_1 , buf_splitterG25ton193n281_n281_4 , 0 , buf_splitterG25ton193n281_n281_5 );
buf_AQFP buf_splitterG25ton193n281_n281_6_( clk_2 , buf_splitterG25ton193n281_n281_5 , 0 , buf_splitterG25ton193n281_n281_6 );
buf_AQFP buf_splitterG25ton193n281_n281_7_( clk_3 , buf_splitterG25ton193n281_n281_6 , 0 , buf_splitterG25ton193n281_n281_7 );
buf_AQFP buf_splitterG25ton193n281_n281_8_( clk_5 , buf_splitterG25ton193n281_n281_7 , 0 , buf_splitterG25ton193n281_n281_8 );
buf_AQFP buf_splitterG25ton193n281_n281_9_( clk_7 , buf_splitterG25ton193n281_n281_8 , 0 , buf_splitterG25ton193n281_n281_9 );
buf_AQFP buf_splitterG26ton100n320_n320_1_( clk_3 , splitterG26ton100n320 , 0 , buf_splitterG26ton100n320_n320_1 );
buf_AQFP buf_splitterG26ton100n320_n320_2_( clk_5 , buf_splitterG26ton100n320_n320_1 , 0 , buf_splitterG26ton100n320_n320_2 );
buf_AQFP buf_splitterG26ton100n320_n320_3_( clk_6 , buf_splitterG26ton100n320_n320_2 , 0 , buf_splitterG26ton100n320_n320_3 );
buf_AQFP buf_splitterG26ton100n320_n320_4_( clk_8 , buf_splitterG26ton100n320_n320_3 , 0 , buf_splitterG26ton100n320_n320_4 );
buf_AQFP buf_splitterG26ton100n320_n320_5_( clk_2 , buf_splitterG26ton100n320_n320_4 , 0 , buf_splitterG26ton100n320_n320_5 );
buf_AQFP buf_splitterG26ton100n320_n320_6_( clk_4 , buf_splitterG26ton100n320_n320_5 , 0 , buf_splitterG26ton100n320_n320_6 );
buf_AQFP buf_splitterG26ton100n320_n320_7_( clk_6 , buf_splitterG26ton100n320_n320_6 , 0 , buf_splitterG26ton100n320_n320_7 );
buf_AQFP buf_splitterG26ton100n320_n320_8_( clk_8 , buf_splitterG26ton100n320_n320_7 , 0 , buf_splitterG26ton100n320_n320_8 );
buf_AQFP buf_splitterG27ton153n287_n287_1_( clk_3 , splitterG27ton153n287 , 0 , buf_splitterG27ton153n287_n287_1 );
buf_AQFP buf_splitterG28ton173n291_n291_1_( clk_3 , splitterG28ton173n291 , 0 , buf_splitterG28ton173n291_n291_1 );
buf_AQFP buf_splitterfromG29_n199_1_( clk_5 , splitterfromG29 , 0 , buf_splitterfromG29_n199_1 );
buf_AQFP buf_splitterG3ton156n46_n213_1_( clk_4 , splitterG3ton156n46 , 0 , buf_splitterG3ton156n46_n213_1 );
buf_AQFP buf_splitterG3ton156n46_n213_2_( clk_6 , buf_splitterG3ton156n46_n213_1 , 0 , buf_splitterG3ton156n46_n213_2 );
buf_AQFP buf_splitterG3ton156n46_n213_3_( clk_8 , buf_splitterG3ton156n46_n213_2 , 0 , buf_splitterG3ton156n46_n213_3 );
buf_AQFP buf_splitterG3ton156n46_n213_4_( clk_2 , buf_splitterG3ton156n46_n213_3 , 0 , buf_splitterG3ton156n46_n213_4 );
buf_AQFP buf_splitterG3ton156n46_n213_5_( clk_4 , buf_splitterG3ton156n46_n213_4 , 0 , buf_splitterG3ton156n46_n213_5 );
buf_AQFP buf_splitterG3ton156n46_n213_6_( clk_5 , buf_splitterG3ton156n46_n213_5 , 0 , buf_splitterG3ton156n46_n213_6 );
buf_AQFP buf_splitterG3ton156n46_n213_7_( clk_6 , buf_splitterG3ton156n46_n213_6 , 0 , buf_splitterG3ton156n46_n213_7 );
buf_AQFP buf_splitterG3ton156n46_n213_8_( clk_8 , buf_splitterG3ton156n46_n213_7 , 0 , buf_splitterG3ton156n46_n213_8 );
buf_AQFP buf_splitterG3ton156n46_n213_9_( clk_2 , buf_splitterG3ton156n46_n213_8 , 0 , buf_splitterG3ton156n46_n213_9 );
buf_AQFP buf_splitterG3ton156n46_n213_10_( clk_4 , buf_splitterG3ton156n46_n213_9 , 0 , buf_splitterG3ton156n46_n213_10 );
buf_AQFP buf_splitterG3ton156n46_n213_11_( clk_6 , buf_splitterG3ton156n46_n213_10 , 0 , buf_splitterG3ton156n46_n213_11 );
buf_AQFP buf_splitterG3ton156n46_n213_12_( clk_8 , buf_splitterG3ton156n46_n213_11 , 0 , buf_splitterG3ton156n46_n213_12 );
buf_AQFP buf_splitterG3ton156n46_n213_13_( clk_2 , buf_splitterG3ton156n46_n213_12 , 0 , buf_splitterG3ton156n46_n213_13 );
buf_AQFP buf_splitterG3ton156n46_n213_14_( clk_4 , buf_splitterG3ton156n46_n213_13 , 0 , buf_splitterG3ton156n46_n213_14 );
buf_AQFP buf_splitterG3ton156n46_n213_15_( clk_6 , buf_splitterG3ton156n46_n213_14 , 0 , buf_splitterG3ton156n46_n213_15 );
buf_AQFP buf_splitterG3ton214n46_n214_1_( clk_5 , splitterG3ton214n46 , 0 , buf_splitterG3ton214n46_n214_1 );
buf_AQFP buf_splitterG3ton214n46_n214_2_( clk_7 , buf_splitterG3ton214n46_n214_1 , 0 , buf_splitterG3ton214n46_n214_2 );
buf_AQFP buf_splitterG3ton214n46_n214_3_( clk_1 , buf_splitterG3ton214n46_n214_2 , 0 , buf_splitterG3ton214n46_n214_3 );
buf_AQFP buf_splitterG3ton214n46_n214_4_( clk_3 , buf_splitterG3ton214n46_n214_3 , 0 , buf_splitterG3ton214n46_n214_4 );
buf_AQFP buf_splitterG3ton214n46_n214_5_( clk_5 , buf_splitterG3ton214n46_n214_4 , 0 , buf_splitterG3ton214n46_n214_5 );
buf_AQFP buf_splitterG3ton214n46_n214_6_( clk_7 , buf_splitterG3ton214n46_n214_5 , 0 , buf_splitterG3ton214n46_n214_6 );
buf_AQFP buf_splitterG3ton214n46_n214_7_( clk_1 , buf_splitterG3ton214n46_n214_6 , 0 , buf_splitterG3ton214n46_n214_7 );
buf_AQFP buf_splitterG3ton214n46_n214_8_( clk_3 , buf_splitterG3ton214n46_n214_7 , 0 , buf_splitterG3ton214n46_n214_8 );
buf_AQFP buf_splitterG3ton214n46_n214_9_( clk_5 , buf_splitterG3ton214n46_n214_8 , 0 , buf_splitterG3ton214n46_n214_9 );
buf_AQFP buf_splitterG3ton214n46_n214_10_( clk_7 , buf_splitterG3ton214n46_n214_9 , 0 , buf_splitterG3ton214n46_n214_10 );
buf_AQFP buf_splitterG3ton214n46_n214_11_( clk_1 , buf_splitterG3ton214n46_n214_10 , 0 , buf_splitterG3ton214n46_n214_11 );
buf_AQFP buf_splitterG3ton214n46_n214_12_( clk_3 , buf_splitterG3ton214n46_n214_11 , 0 , buf_splitterG3ton214n46_n214_12 );
buf_AQFP buf_splitterG3ton214n46_n214_13_( clk_5 , buf_splitterG3ton214n46_n214_12 , 0 , buf_splitterG3ton214n46_n214_13 );
buf_AQFP buf_splitterfromG30_n312_1_( clk_5 , splitterfromG30 , 0 , buf_splitterfromG30_n312_1 );
buf_AQFP buf_splitterG31ton126n127_n126_1_( clk_6 , splitterG31ton126n127 , 0 , buf_splitterG31ton126n127_n126_1 );
buf_AQFP buf_splitterG31ton126n127_n126_2_( clk_8 , buf_splitterG31ton126n127_n126_1 , 0 , buf_splitterG31ton126n127_n126_2 );
buf_AQFP buf_splitterG31ton152n201_n152_1_( clk_6 , splitterG31ton152n201 , 0 , buf_splitterG31ton152n201_n152_1 );
buf_AQFP buf_splitterG31ton152n201_n152_2_( clk_7 , buf_splitterG31ton152n201_n152_1 , 0 , buf_splitterG31ton152n201_n152_2 );
buf_AQFP buf_splitterG31ton152n201_n172_1_( clk_7 , splitterG31ton152n201 , 0 , buf_splitterG31ton152n201_n172_1 );
buf_AQFP buf_splitterG31ton152n201_n192_1_( clk_6 , splitterG31ton152n201 , 0 , buf_splitterG31ton152n201_n192_1 );
buf_AQFP buf_splitterG31ton152n201_n192_2_( clk_8 , buf_splitterG31ton152n201_n192_1 , 0 , buf_splitterG31ton152n201_n192_2 );
buf_AQFP buf_splitterG31ton276n291_n276_1_( clk_5 , splitterG31ton276n291 , 0 , buf_splitterG31ton276n291_n276_1 );
buf_AQFP buf_splitterG31ton276n291_n276_2_( clk_6 , buf_splitterG31ton276n291_n276_1 , 0 , buf_splitterG31ton276n291_n276_2 );
buf_AQFP buf_splitterG31ton276n291_n276_3_( clk_8 , buf_splitterG31ton276n291_n276_2 , 0 , buf_splitterG31ton276n291_n276_3 );
buf_AQFP buf_splitterG31ton276n291_n276_4_( clk_2 , buf_splitterG31ton276n291_n276_3 , 0 , buf_splitterG31ton276n291_n276_4 );
buf_AQFP buf_splitterG31ton276n291_n276_5_( clk_4 , buf_splitterG31ton276n291_n276_4 , 0 , buf_splitterG31ton276n291_n276_5 );
buf_AQFP buf_splitterG31ton276n291_n276_6_( clk_6 , buf_splitterG31ton276n291_n276_5 , 0 , buf_splitterG31ton276n291_n276_6 );
buf_AQFP buf_splitterG31ton276n291_n276_7_( clk_7 , buf_splitterG31ton276n291_n276_6 , 0 , buf_splitterG31ton276n291_n276_7 );
buf_AQFP buf_splitterG31ton276n291_n276_8_( clk_1 , buf_splitterG31ton276n291_n276_7 , 0 , buf_splitterG31ton276n291_n276_8 );
buf_AQFP buf_splitterG31ton276n291_n282_1_( clk_5 , splitterG31ton276n291 , 0 , buf_splitterG31ton276n291_n282_1 );
buf_AQFP buf_splitterG31ton276n291_n282_2_( clk_7 , buf_splitterG31ton276n291_n282_1 , 0 , buf_splitterG31ton276n291_n282_2 );
buf_AQFP buf_splitterG31ton276n291_n282_3_( clk_1 , buf_splitterG31ton276n291_n282_2 , 0 , buf_splitterG31ton276n291_n282_3 );
buf_AQFP buf_splitterG31ton276n291_n282_4_( clk_2 , buf_splitterG31ton276n291_n282_3 , 0 , buf_splitterG31ton276n291_n282_4 );
buf_AQFP buf_splitterG31ton276n291_n282_5_( clk_4 , buf_splitterG31ton276n291_n282_4 , 0 , buf_splitterG31ton276n291_n282_5 );
buf_AQFP buf_splitterG31ton276n291_n282_6_( clk_6 , buf_splitterG31ton276n291_n282_5 , 0 , buf_splitterG31ton276n291_n282_6 );
buf_AQFP buf_splitterG31ton276n291_n282_7_( clk_7 , buf_splitterG31ton276n291_n282_6 , 0 , buf_splitterG31ton276n291_n282_7 );
buf_AQFP buf_splitterG31ton276n291_n282_8_( clk_1 , buf_splitterG31ton276n291_n282_7 , 0 , buf_splitterG31ton276n291_n282_8 );
buf_AQFP buf_splitterG31ton295n99_n295_1_( clk_4 , splitterG31ton295n99 , 0 , buf_splitterG31ton295n99_n295_1 );
buf_AQFP buf_splitterG31ton295n99_n295_2_( clk_6 , buf_splitterG31ton295n99_n295_1 , 0 , buf_splitterG31ton295n99_n295_2 );
buf_AQFP buf_splitterG31ton295n99_n295_3_( clk_8 , buf_splitterG31ton295n99_n295_2 , 0 , buf_splitterG31ton295n99_n295_3 );
buf_AQFP buf_splitterG31ton295n99_n295_4_( clk_2 , buf_splitterG31ton295n99_n295_3 , 0 , buf_splitterG31ton295n99_n295_4 );
buf_AQFP buf_splitterG31ton295n99_n295_5_( clk_4 , buf_splitterG31ton295n99_n295_4 , 0 , buf_splitterG31ton295n99_n295_5 );
buf_AQFP buf_splitterG31ton295n99_n73_1_( clk_3 , splitterG31ton295n99 , 0 , buf_splitterG31ton295n99_n73_1 );
buf_AQFP buf_splitterG31ton295n99_n73_2_( clk_5 , buf_splitterG31ton295n99_n73_1 , 0 , buf_splitterG31ton295n99_n73_2 );
buf_AQFP buf_splitterG31ton295n99_n73_3_( clk_6 , buf_splitterG31ton295n99_n73_2 , 0 , buf_splitterG31ton295n99_n73_3 );
buf_AQFP buf_splitterG31ton295n99_n73_4_( clk_7 , buf_splitterG31ton295n99_n73_3 , 0 , buf_splitterG31ton295n99_n73_4 );
buf_AQFP buf_splitterG31ton295n99_n73_5_( clk_1 , buf_splitterG31ton295n99_n73_4 , 0 , buf_splitterG31ton295n99_n73_5 );
buf_AQFP buf_splitterG31ton295n99_n99_1_( clk_4 , splitterG31ton295n99 , 0 , buf_splitterG31ton295n99_n99_1 );
buf_AQFP buf_splitterG31ton295n99_n99_2_( clk_5 , buf_splitterG31ton295n99_n99_1 , 0 , buf_splitterG31ton295n99_n99_2 );
buf_AQFP buf_splitterG31ton295n99_n99_3_( clk_7 , buf_splitterG31ton295n99_n99_2 , 0 , buf_splitterG31ton295n99_n99_3 );
buf_AQFP buf_splitterfromG32_n268_1_( clk_7 , splitterfromG32 , 0 , buf_splitterfromG32_n268_1 );
buf_AQFP buf_splitterfromG32_n268_2_( clk_1 , buf_splitterfromG32_n268_1 , 0 , buf_splitterfromG32_n268_2 );
buf_AQFP buf_splitterfromG32_n268_3_( clk_3 , buf_splitterfromG32_n268_2 , 0 , buf_splitterfromG32_n268_3 );
buf_AQFP buf_splitterfromG32_n268_4_( clk_5 , buf_splitterfromG32_n268_3 , 0 , buf_splitterfromG32_n268_4 );
buf_AQFP buf_splitterfromG32_n268_5_( clk_7 , buf_splitterfromG32_n268_4 , 0 , buf_splitterfromG32_n268_5 );
buf_AQFP buf_splitterfromG32_n268_6_( clk_1 , buf_splitterfromG32_n268_5 , 0 , buf_splitterfromG32_n268_6 );
buf_AQFP buf_splitterfromG32_n268_7_( clk_3 , buf_splitterfromG32_n268_6 , 0 , buf_splitterfromG32_n268_7 );
buf_AQFP buf_splitterfromG32_n268_8_( clk_5 , buf_splitterfromG32_n268_7 , 0 , buf_splitterfromG32_n268_8 );
buf_AQFP buf_splitterfromG32_n268_9_( clk_7 , buf_splitterfromG32_n268_8 , 0 , buf_splitterfromG32_n268_9 );
buf_AQFP buf_splitterfromG32_n268_10_( clk_1 , buf_splitterfromG32_n268_9 , 0 , buf_splitterfromG32_n268_10 );
buf_AQFP buf_splitterfromG32_n268_11_( clk_3 , buf_splitterfromG32_n268_10 , 0 , buf_splitterfromG32_n268_11 );
buf_AQFP buf_splitterfromG32_n268_12_( clk_5 , buf_splitterfromG32_n268_11 , 0 , buf_splitterfromG32_n268_12 );
buf_AQFP buf_splitterfromG32_n268_13_( clk_7 , buf_splitterfromG32_n268_12 , 0 , buf_splitterfromG32_n268_13 );
buf_AQFP buf_splitterfromG32_n268_14_( clk_8 , buf_splitterfromG32_n268_13 , 0 , buf_splitterfromG32_n268_14 );
buf_AQFP buf_splitterG33ton109n88_n179_1_( clk_3 , splitterG33ton109n88 , 0 , buf_splitterG33ton109n88_n179_1 );
buf_AQFP buf_splitterG33ton199n273_n203_1_( clk_5 , splitterG33ton199n273 , 0 , buf_splitterG33ton199n273_n203_1 );
buf_AQFP buf_splitterG33ton199n273_n273_1_( clk_6 , splitterG33ton199n273 , 0 , buf_splitterG33ton199n273_n273_1 );
buf_AQFP buf_splitterG33ton199n273_n273_2_( clk_8 , buf_splitterG33ton199n273_n273_1 , 0 , buf_splitterG33ton199n273_n273_2 );
buf_AQFP buf_splitterG33ton199n273_n273_3_( clk_2 , buf_splitterG33ton199n273_n273_2 , 0 , buf_splitterG33ton199n273_n273_3 );
buf_AQFP buf_splitterG33ton199n273_n273_4_( clk_4 , buf_splitterG33ton199n273_n273_3 , 0 , buf_splitterG33ton199n273_n273_4 );
buf_AQFP buf_splitterG33ton199n273_n273_5_( clk_6 , buf_splitterG33ton199n273_n273_4 , 0 , buf_splitterG33ton199n273_n273_5 );
buf_AQFP buf_splitterG33ton199n273_n273_6_( clk_8 , buf_splitterG33ton199n273_n273_5 , 0 , buf_splitterG33ton199n273_n273_6 );
buf_AQFP buf_splitterG33ton199n273_n273_7_( clk_2 , buf_splitterG33ton199n273_n273_6 , 0 , buf_splitterG33ton199n273_n273_7 );
buf_AQFP buf_splitterG33ton199n273_n273_8_( clk_4 , buf_splitterG33ton199n273_n273_7 , 0 , buf_splitterG33ton199n273_n273_8 );
buf_AQFP buf_splitterG33ton199n273_n273_9_( clk_6 , buf_splitterG33ton199n273_n273_8 , 0 , buf_splitterG33ton199n273_n273_9 );
buf_AQFP buf_splitterG33ton199n273_n273_10_( clk_8 , buf_splitterG33ton199n273_n273_9 , 0 , buf_splitterG33ton199n273_n273_10 );
buf_AQFP buf_splitterG33ton199n273_n273_11_( clk_2 , buf_splitterG33ton199n273_n273_10 , 0 , buf_splitterG33ton199n273_n273_11 );
buf_AQFP buf_splitterG33ton304n88_n304_1_( clk_5 , splitterG33ton304n88 , 0 , buf_splitterG33ton304n88_n304_1 );
buf_AQFP buf_splitterG33ton304n88_n304_2_( clk_7 , buf_splitterG33ton304n88_n304_1 , 0 , buf_splitterG33ton304n88_n304_2 );
buf_AQFP buf_splitterG33ton304n88_n304_3_( clk_1 , buf_splitterG33ton304n88_n304_2 , 0 , buf_splitterG33ton304n88_n304_3 );
buf_AQFP buf_splitterG33ton304n88_n304_4_( clk_3 , buf_splitterG33ton304n88_n304_3 , 0 , buf_splitterG33ton304n88_n304_4 );
buf_AQFP buf_splitterG33ton304n88_n304_5_( clk_5 , buf_splitterG33ton304n88_n304_4 , 0 , buf_splitterG33ton304n88_n304_5 );
buf_AQFP buf_splitterG33ton304n88_n304_6_( clk_7 , buf_splitterG33ton304n88_n304_5 , 0 , buf_splitterG33ton304n88_n304_6 );
buf_AQFP buf_splitterG33ton304n88_n304_7_( clk_1 , buf_splitterG33ton304n88_n304_6 , 0 , buf_splitterG33ton304n88_n304_7 );
buf_AQFP buf_splitterG33ton304n88_n304_8_( clk_3 , buf_splitterG33ton304n88_n304_7 , 0 , buf_splitterG33ton304n88_n304_8 );
buf_AQFP buf_splitterG33ton304n88_n304_9_( clk_5 , buf_splitterG33ton304n88_n304_8 , 0 , buf_splitterG33ton304n88_n304_9 );
buf_AQFP buf_splitterG33ton304n88_n304_10_( clk_7 , buf_splitterG33ton304n88_n304_9 , 0 , buf_splitterG33ton304n88_n304_10 );
buf_AQFP buf_splitterG33ton304n88_n304_11_( clk_1 , buf_splitterG33ton304n88_n304_10 , 0 , buf_splitterG33ton304n88_n304_11 );
buf_AQFP buf_splitterG33ton304n88_n304_12_( clk_3 , buf_splitterG33ton304n88_n304_11 , 0 , buf_splitterG33ton304n88_n304_12 );
buf_AQFP buf_splitterG33ton304n88_n304_13_( clk_5 , buf_splitterG33ton304n88_n304_12 , 0 , buf_splitterG33ton304n88_n304_13 );
buf_AQFP buf_splitterG33ton304n88_n304_14_( clk_7 , buf_splitterG33ton304n88_n304_13 , 0 , buf_splitterG33ton304n88_n304_14 );
buf_AQFP buf_splitterG33ton304n88_n316_1_( clk_5 , splitterG33ton304n88 , 0 , buf_splitterG33ton304n88_n316_1 );
buf_AQFP buf_splitterG33ton304n88_n316_2_( clk_7 , buf_splitterG33ton304n88_n316_1 , 0 , buf_splitterG33ton304n88_n316_2 );
buf_AQFP buf_splitterG33ton304n88_n316_3_( clk_1 , buf_splitterG33ton304n88_n316_2 , 0 , buf_splitterG33ton304n88_n316_3 );
buf_AQFP buf_splitterG33ton304n88_n316_4_( clk_3 , buf_splitterG33ton304n88_n316_3 , 0 , buf_splitterG33ton304n88_n316_4 );
buf_AQFP buf_splitterG33ton304n88_n316_5_( clk_5 , buf_splitterG33ton304n88_n316_4 , 0 , buf_splitterG33ton304n88_n316_5 );
buf_AQFP buf_splitterG33ton304n88_n316_6_( clk_7 , buf_splitterG33ton304n88_n316_5 , 0 , buf_splitterG33ton304n88_n316_6 );
buf_AQFP buf_splitterG33ton304n88_n316_7_( clk_1 , buf_splitterG33ton304n88_n316_6 , 0 , buf_splitterG33ton304n88_n316_7 );
buf_AQFP buf_splitterG33ton304n88_n316_8_( clk_3 , buf_splitterG33ton304n88_n316_7 , 0 , buf_splitterG33ton304n88_n316_8 );
buf_AQFP buf_splitterG33ton304n88_n316_9_( clk_5 , buf_splitterG33ton304n88_n316_8 , 0 , buf_splitterG33ton304n88_n316_9 );
buf_AQFP buf_splitterG33ton304n88_n316_10_( clk_7 , buf_splitterG33ton304n88_n316_9 , 0 , buf_splitterG33ton304n88_n316_10 );
buf_AQFP buf_splitterG33ton304n88_n316_11_( clk_8 , buf_splitterG33ton304n88_n316_10 , 0 , buf_splitterG33ton304n88_n316_11 );
buf_AQFP buf_splitterG33ton304n88_n316_12_( clk_1 , buf_splitterG33ton304n88_n316_11 , 0 , buf_splitterG33ton304n88_n316_12 );
buf_AQFP buf_splitterG33ton304n88_n316_13_( clk_3 , buf_splitterG33ton304n88_n316_12 , 0 , buf_splitterG33ton304n88_n316_13 );
buf_AQFP buf_splitterG33ton304n88_n316_14_( clk_5 , buf_splitterG33ton304n88_n316_13 , 0 , buf_splitterG33ton304n88_n316_14 );
buf_AQFP buf_splitterG33ton304n88_n316_15_( clk_6 , buf_splitterG33ton304n88_n316_14 , 0 , buf_splitterG33ton304n88_n316_15 );
buf_AQFP buf_splitterG33ton304n88_n316_16_( clk_7 , buf_splitterG33ton304n88_n316_15 , 0 , buf_splitterG33ton304n88_n316_16 );
buf_AQFP buf_splitterG4ton216n43_n216_1_( clk_8 , splitterG4ton216n43 , 0 , buf_splitterG4ton216n43_n216_1 );
buf_AQFP buf_splitterG4ton216n43_n216_2_( clk_2 , buf_splitterG4ton216n43_n216_1 , 0 , buf_splitterG4ton216n43_n216_2 );
buf_AQFP buf_splitterG4ton216n43_n216_3_( clk_4 , buf_splitterG4ton216n43_n216_2 , 0 , buf_splitterG4ton216n43_n216_3 );
buf_AQFP buf_splitterG4ton216n43_n216_4_( clk_6 , buf_splitterG4ton216n43_n216_3 , 0 , buf_splitterG4ton216n43_n216_4 );
buf_AQFP buf_splitterG4ton216n43_n216_5_( clk_8 , buf_splitterG4ton216n43_n216_4 , 0 , buf_splitterG4ton216n43_n216_5 );
buf_AQFP buf_splitterG4ton216n43_n216_6_( clk_2 , buf_splitterG4ton216n43_n216_5 , 0 , buf_splitterG4ton216n43_n216_6 );
buf_AQFP buf_splitterG4ton216n43_n216_7_( clk_4 , buf_splitterG4ton216n43_n216_6 , 0 , buf_splitterG4ton216n43_n216_7 );
buf_AQFP buf_splitterG4ton216n43_n216_8_( clk_6 , buf_splitterG4ton216n43_n216_7 , 0 , buf_splitterG4ton216n43_n216_8 );
buf_AQFP buf_splitterG4ton216n43_n216_9_( clk_8 , buf_splitterG4ton216n43_n216_8 , 0 , buf_splitterG4ton216n43_n216_9 );
buf_AQFP buf_splitterG4ton216n43_n216_10_( clk_1 , buf_splitterG4ton216n43_n216_9 , 0 , buf_splitterG4ton216n43_n216_10 );
buf_AQFP buf_splitterG4ton216n43_n216_11_( clk_3 , buf_splitterG4ton216n43_n216_10 , 0 , buf_splitterG4ton216n43_n216_11 );
buf_AQFP buf_splitterG4ton216n43_n216_12_( clk_4 , buf_splitterG4ton216n43_n216_11 , 0 , buf_splitterG4ton216n43_n216_12 );
buf_AQFP buf_splitterG4ton216n43_n216_13_( clk_6 , buf_splitterG4ton216n43_n216_12 , 0 , buf_splitterG4ton216n43_n216_13 );
buf_AQFP buf_splitterG4ton216n43_n217_1_( clk_8 , splitterG4ton216n43 , 0 , buf_splitterG4ton216n43_n217_1 );
buf_AQFP buf_splitterG4ton216n43_n217_2_( clk_2 , buf_splitterG4ton216n43_n217_1 , 0 , buf_splitterG4ton216n43_n217_2 );
buf_AQFP buf_splitterG4ton216n43_n217_3_( clk_4 , buf_splitterG4ton216n43_n217_2 , 0 , buf_splitterG4ton216n43_n217_3 );
buf_AQFP buf_splitterG4ton216n43_n217_4_( clk_6 , buf_splitterG4ton216n43_n217_3 , 0 , buf_splitterG4ton216n43_n217_4 );
buf_AQFP buf_splitterG4ton216n43_n217_5_( clk_8 , buf_splitterG4ton216n43_n217_4 , 0 , buf_splitterG4ton216n43_n217_5 );
buf_AQFP buf_splitterG4ton216n43_n217_6_( clk_2 , buf_splitterG4ton216n43_n217_5 , 0 , buf_splitterG4ton216n43_n217_6 );
buf_AQFP buf_splitterG4ton216n43_n217_7_( clk_3 , buf_splitterG4ton216n43_n217_6 , 0 , buf_splitterG4ton216n43_n217_7 );
buf_AQFP buf_splitterG4ton216n43_n217_8_( clk_5 , buf_splitterG4ton216n43_n217_7 , 0 , buf_splitterG4ton216n43_n217_8 );
buf_AQFP buf_splitterG4ton216n43_n217_9_( clk_7 , buf_splitterG4ton216n43_n217_8 , 0 , buf_splitterG4ton216n43_n217_9 );
buf_AQFP buf_splitterG4ton216n43_n217_10_( clk_1 , buf_splitterG4ton216n43_n217_9 , 0 , buf_splitterG4ton216n43_n217_10 );
buf_AQFP buf_splitterG4ton216n43_n217_11_( clk_3 , buf_splitterG4ton216n43_n217_10 , 0 , buf_splitterG4ton216n43_n217_11 );
buf_AQFP buf_splitterG4ton216n43_n217_12_( clk_5 , buf_splitterG4ton216n43_n217_11 , 0 , buf_splitterG4ton216n43_n217_12 );
buf_AQFP buf_splitterG5ton143n40_n236_1_( clk_4 , splitterG5ton143n40 , 0 , buf_splitterG5ton143n40_n236_1 );
buf_AQFP buf_splitterG5ton143n40_n236_2_( clk_6 , buf_splitterG5ton143n40_n236_1 , 0 , buf_splitterG5ton143n40_n236_2 );
buf_AQFP buf_splitterG5ton143n40_n236_3_( clk_8 , buf_splitterG5ton143n40_n236_2 , 0 , buf_splitterG5ton143n40_n236_3 );
buf_AQFP buf_splitterG5ton143n40_n236_4_( clk_2 , buf_splitterG5ton143n40_n236_3 , 0 , buf_splitterG5ton143n40_n236_4 );
buf_AQFP buf_splitterG5ton143n40_n236_5_( clk_4 , buf_splitterG5ton143n40_n236_4 , 0 , buf_splitterG5ton143n40_n236_5 );
buf_AQFP buf_splitterG5ton143n40_n236_6_( clk_6 , buf_splitterG5ton143n40_n236_5 , 0 , buf_splitterG5ton143n40_n236_6 );
buf_AQFP buf_splitterG5ton143n40_n236_7_( clk_8 , buf_splitterG5ton143n40_n236_6 , 0 , buf_splitterG5ton143n40_n236_7 );
buf_AQFP buf_splitterG5ton143n40_n236_8_( clk_2 , buf_splitterG5ton143n40_n236_7 , 0 , buf_splitterG5ton143n40_n236_8 );
buf_AQFP buf_splitterG5ton143n40_n236_9_( clk_4 , buf_splitterG5ton143n40_n236_8 , 0 , buf_splitterG5ton143n40_n236_9 );
buf_AQFP buf_splitterG5ton143n40_n236_10_( clk_6 , buf_splitterG5ton143n40_n236_9 , 0 , buf_splitterG5ton143n40_n236_10 );
buf_AQFP buf_splitterG5ton143n40_n236_11_( clk_8 , buf_splitterG5ton143n40_n236_10 , 0 , buf_splitterG5ton143n40_n236_11 );
buf_AQFP buf_splitterG5ton143n40_n236_12_( clk_2 , buf_splitterG5ton143n40_n236_11 , 0 , buf_splitterG5ton143n40_n236_12 );
buf_AQFP buf_splitterG5ton143n40_n236_13_( clk_4 , buf_splitterG5ton143n40_n236_12 , 0 , buf_splitterG5ton143n40_n236_13 );
buf_AQFP buf_splitterG5ton237n40_n237_1_( clk_1 , splitterG5ton237n40 , 0 , buf_splitterG5ton237n40_n237_1 );
buf_AQFP buf_splitterG5ton237n40_n237_2_( clk_3 , buf_splitterG5ton237n40_n237_1 , 0 , buf_splitterG5ton237n40_n237_2 );
buf_AQFP buf_splitterG5ton237n40_n237_3_( clk_5 , buf_splitterG5ton237n40_n237_2 , 0 , buf_splitterG5ton237n40_n237_3 );
buf_AQFP buf_splitterG5ton237n40_n237_4_( clk_7 , buf_splitterG5ton237n40_n237_3 , 0 , buf_splitterG5ton237n40_n237_4 );
buf_AQFP buf_splitterG5ton237n40_n237_5_( clk_1 , buf_splitterG5ton237n40_n237_4 , 0 , buf_splitterG5ton237n40_n237_5 );
buf_AQFP buf_splitterG5ton237n40_n237_6_( clk_3 , buf_splitterG5ton237n40_n237_5 , 0 , buf_splitterG5ton237n40_n237_6 );
buf_AQFP buf_splitterG5ton237n40_n237_7_( clk_5 , buf_splitterG5ton237n40_n237_6 , 0 , buf_splitterG5ton237n40_n237_7 );
buf_AQFP buf_splitterG5ton237n40_n237_8_( clk_7 , buf_splitterG5ton237n40_n237_7 , 0 , buf_splitterG5ton237n40_n237_8 );
buf_AQFP buf_splitterG5ton237n40_n237_9_( clk_1 , buf_splitterG5ton237n40_n237_8 , 0 , buf_splitterG5ton237n40_n237_9 );
buf_AQFP buf_splitterG5ton237n40_n237_10_( clk_2 , buf_splitterG5ton237n40_n237_9 , 0 , buf_splitterG5ton237n40_n237_10 );
buf_AQFP buf_splitterG5ton237n40_n237_11_( clk_4 , buf_splitterG5ton237n40_n237_10 , 0 , buf_splitterG5ton237n40_n237_11 );
buf_AQFP buf_splitterG6ton156n37_n239_1_( clk_5 , splitterG6ton156n37 , 0 , buf_splitterG6ton156n37_n239_1 );
buf_AQFP buf_splitterG6ton156n37_n239_2_( clk_7 , buf_splitterG6ton156n37_n239_1 , 0 , buf_splitterG6ton156n37_n239_2 );
buf_AQFP buf_splitterG6ton156n37_n239_3_( clk_1 , buf_splitterG6ton156n37_n239_2 , 0 , buf_splitterG6ton156n37_n239_3 );
buf_AQFP buf_splitterG6ton156n37_n239_4_( clk_3 , buf_splitterG6ton156n37_n239_3 , 0 , buf_splitterG6ton156n37_n239_4 );
buf_AQFP buf_splitterG6ton156n37_n239_5_( clk_5 , buf_splitterG6ton156n37_n239_4 , 0 , buf_splitterG6ton156n37_n239_5 );
buf_AQFP buf_splitterG6ton156n37_n239_6_( clk_7 , buf_splitterG6ton156n37_n239_5 , 0 , buf_splitterG6ton156n37_n239_6 );
buf_AQFP buf_splitterG6ton156n37_n239_7_( clk_1 , buf_splitterG6ton156n37_n239_6 , 0 , buf_splitterG6ton156n37_n239_7 );
buf_AQFP buf_splitterG6ton156n37_n239_8_( clk_2 , buf_splitterG6ton156n37_n239_7 , 0 , buf_splitterG6ton156n37_n239_8 );
buf_AQFP buf_splitterG6ton156n37_n239_9_( clk_4 , buf_splitterG6ton156n37_n239_8 , 0 , buf_splitterG6ton156n37_n239_9 );
buf_AQFP buf_splitterG6ton156n37_n239_10_( clk_6 , buf_splitterG6ton156n37_n239_9 , 0 , buf_splitterG6ton156n37_n239_10 );
buf_AQFP buf_splitterG6ton156n37_n239_11_( clk_8 , buf_splitterG6ton156n37_n239_10 , 0 , buf_splitterG6ton156n37_n239_11 );
buf_AQFP buf_splitterG6ton156n37_n239_12_( clk_2 , buf_splitterG6ton156n37_n239_11 , 0 , buf_splitterG6ton156n37_n239_12 );
buf_AQFP buf_splitterG6ton156n37_n239_13_( clk_4 , buf_splitterG6ton156n37_n239_12 , 0 , buf_splitterG6ton156n37_n239_13 );
buf_AQFP buf_splitterG6ton156n37_n239_14_( clk_6 , buf_splitterG6ton156n37_n239_13 , 0 , buf_splitterG6ton156n37_n239_14 );
buf_AQFP buf_splitterG6ton240n37_n240_1_( clk_6 , splitterG6ton240n37 , 0 , buf_splitterG6ton240n37_n240_1 );
buf_AQFP buf_splitterG6ton240n37_n240_2_( clk_8 , buf_splitterG6ton240n37_n240_1 , 0 , buf_splitterG6ton240n37_n240_2 );
buf_AQFP buf_splitterG6ton240n37_n240_3_( clk_2 , buf_splitterG6ton240n37_n240_2 , 0 , buf_splitterG6ton240n37_n240_3 );
buf_AQFP buf_splitterG6ton240n37_n240_4_( clk_4 , buf_splitterG6ton240n37_n240_3 , 0 , buf_splitterG6ton240n37_n240_4 );
buf_AQFP buf_splitterG6ton240n37_n240_5_( clk_6 , buf_splitterG6ton240n37_n240_4 , 0 , buf_splitterG6ton240n37_n240_5 );
buf_AQFP buf_splitterG6ton240n37_n240_6_( clk_8 , buf_splitterG6ton240n37_n240_5 , 0 , buf_splitterG6ton240n37_n240_6 );
buf_AQFP buf_splitterG6ton240n37_n240_7_( clk_2 , buf_splitterG6ton240n37_n240_6 , 0 , buf_splitterG6ton240n37_n240_7 );
buf_AQFP buf_splitterG6ton240n37_n240_8_( clk_4 , buf_splitterG6ton240n37_n240_7 , 0 , buf_splitterG6ton240n37_n240_8 );
buf_AQFP buf_splitterG6ton240n37_n240_9_( clk_6 , buf_splitterG6ton240n37_n240_8 , 0 , buf_splitterG6ton240n37_n240_9 );
buf_AQFP buf_splitterG6ton240n37_n240_10_( clk_8 , buf_splitterG6ton240n37_n240_9 , 0 , buf_splitterG6ton240n37_n240_10 );
buf_AQFP buf_splitterG6ton240n37_n240_11_( clk_1 , buf_splitterG6ton240n37_n240_10 , 0 , buf_splitterG6ton240n37_n240_11 );
buf_AQFP buf_splitterG6ton240n37_n240_12_( clk_3 , buf_splitterG6ton240n37_n240_11 , 0 , buf_splitterG6ton240n37_n240_12 );
buf_AQFP buf_splitterG6ton240n37_n240_13_( clk_5 , buf_splitterG6ton240n37_n240_12 , 0 , buf_splitterG6ton240n37_n240_13 );
buf_AQFP buf_splitterG7ton117n37_n242_1_( clk_4 , splitterG7ton117n37 , 0 , buf_splitterG7ton117n37_n242_1 );
buf_AQFP buf_splitterG7ton117n37_n242_2_( clk_6 , buf_splitterG7ton117n37_n242_1 , 0 , buf_splitterG7ton117n37_n242_2 );
buf_AQFP buf_splitterG7ton117n37_n242_3_( clk_8 , buf_splitterG7ton117n37_n242_2 , 0 , buf_splitterG7ton117n37_n242_3 );
buf_AQFP buf_splitterG7ton117n37_n242_4_( clk_2 , buf_splitterG7ton117n37_n242_3 , 0 , buf_splitterG7ton117n37_n242_4 );
buf_AQFP buf_splitterG7ton117n37_n242_5_( clk_4 , buf_splitterG7ton117n37_n242_4 , 0 , buf_splitterG7ton117n37_n242_5 );
buf_AQFP buf_splitterG7ton117n37_n242_6_( clk_6 , buf_splitterG7ton117n37_n242_5 , 0 , buf_splitterG7ton117n37_n242_6 );
buf_AQFP buf_splitterG7ton117n37_n242_7_( clk_8 , buf_splitterG7ton117n37_n242_6 , 0 , buf_splitterG7ton117n37_n242_7 );
buf_AQFP buf_splitterG7ton117n37_n242_8_( clk_2 , buf_splitterG7ton117n37_n242_7 , 0 , buf_splitterG7ton117n37_n242_8 );
buf_AQFP buf_splitterG7ton117n37_n242_9_( clk_4 , buf_splitterG7ton117n37_n242_8 , 0 , buf_splitterG7ton117n37_n242_9 );
buf_AQFP buf_splitterG7ton117n37_n242_10_( clk_6 , buf_splitterG7ton117n37_n242_9 , 0 , buf_splitterG7ton117n37_n242_10 );
buf_AQFP buf_splitterG7ton117n37_n242_11_( clk_8 , buf_splitterG7ton117n37_n242_10 , 0 , buf_splitterG7ton117n37_n242_11 );
buf_AQFP buf_splitterG7ton117n37_n242_12_( clk_2 , buf_splitterG7ton117n37_n242_11 , 0 , buf_splitterG7ton117n37_n242_12 );
buf_AQFP buf_splitterG7ton117n37_n242_13_( clk_4 , buf_splitterG7ton117n37_n242_12 , 0 , buf_splitterG7ton117n37_n242_13 );
buf_AQFP buf_splitterG7ton117n37_n242_14_( clk_6 , buf_splitterG7ton117n37_n242_13 , 0 , buf_splitterG7ton117n37_n242_14 );
buf_AQFP buf_splitterG7ton243n37_n243_1_( clk_6 , splitterG7ton243n37 , 0 , buf_splitterG7ton243n37_n243_1 );
buf_AQFP buf_splitterG7ton243n37_n243_2_( clk_8 , buf_splitterG7ton243n37_n243_1 , 0 , buf_splitterG7ton243n37_n243_2 );
buf_AQFP buf_splitterG7ton243n37_n243_3_( clk_2 , buf_splitterG7ton243n37_n243_2 , 0 , buf_splitterG7ton243n37_n243_3 );
buf_AQFP buf_splitterG7ton243n37_n243_4_( clk_4 , buf_splitterG7ton243n37_n243_3 , 0 , buf_splitterG7ton243n37_n243_4 );
buf_AQFP buf_splitterG7ton243n37_n243_5_( clk_6 , buf_splitterG7ton243n37_n243_4 , 0 , buf_splitterG7ton243n37_n243_5 );
buf_AQFP buf_splitterG7ton243n37_n243_6_( clk_8 , buf_splitterG7ton243n37_n243_5 , 0 , buf_splitterG7ton243n37_n243_6 );
buf_AQFP buf_splitterG7ton243n37_n243_7_( clk_2 , buf_splitterG7ton243n37_n243_6 , 0 , buf_splitterG7ton243n37_n243_7 );
buf_AQFP buf_splitterG7ton243n37_n243_8_( clk_4 , buf_splitterG7ton243n37_n243_7 , 0 , buf_splitterG7ton243n37_n243_8 );
buf_AQFP buf_splitterG7ton243n37_n243_9_( clk_6 , buf_splitterG7ton243n37_n243_8 , 0 , buf_splitterG7ton243n37_n243_9 );
buf_AQFP buf_splitterG7ton243n37_n243_10_( clk_8 , buf_splitterG7ton243n37_n243_9 , 0 , buf_splitterG7ton243n37_n243_10 );
buf_AQFP buf_splitterG7ton243n37_n243_11_( clk_1 , buf_splitterG7ton243n37_n243_10 , 0 , buf_splitterG7ton243n37_n243_11 );
buf_AQFP buf_splitterG7ton243n37_n243_12_( clk_2 , buf_splitterG7ton243n37_n243_11 , 0 , buf_splitterG7ton243n37_n243_12 );
buf_AQFP buf_splitterG7ton243n37_n243_13_( clk_3 , buf_splitterG7ton243n37_n243_12 , 0 , buf_splitterG7ton243n37_n243_13 );
buf_AQFP buf_splitterG7ton243n37_n243_14_( clk_4 , buf_splitterG7ton243n37_n243_13 , 0 , buf_splitterG7ton243n37_n243_14 );
buf_AQFP buf_splitterG7ton243n37_n243_15_( clk_5 , buf_splitterG7ton243n37_n243_14 , 0 , buf_splitterG7ton243n37_n243_15 );
buf_AQFP buf_splitterG8ton245n43_n245_1_( clk_8 , splitterG8ton245n43 , 0 , buf_splitterG8ton245n43_n245_1 );
buf_AQFP buf_splitterG8ton245n43_n245_2_( clk_2 , buf_splitterG8ton245n43_n245_1 , 0 , buf_splitterG8ton245n43_n245_2 );
buf_AQFP buf_splitterG8ton245n43_n245_3_( clk_4 , buf_splitterG8ton245n43_n245_2 , 0 , buf_splitterG8ton245n43_n245_3 );
buf_AQFP buf_splitterG8ton245n43_n245_4_( clk_6 , buf_splitterG8ton245n43_n245_3 , 0 , buf_splitterG8ton245n43_n245_4 );
buf_AQFP buf_splitterG8ton245n43_n245_5_( clk_8 , buf_splitterG8ton245n43_n245_4 , 0 , buf_splitterG8ton245n43_n245_5 );
buf_AQFP buf_splitterG8ton245n43_n245_6_( clk_2 , buf_splitterG8ton245n43_n245_5 , 0 , buf_splitterG8ton245n43_n245_6 );
buf_AQFP buf_splitterG8ton245n43_n245_7_( clk_4 , buf_splitterG8ton245n43_n245_6 , 0 , buf_splitterG8ton245n43_n245_7 );
buf_AQFP buf_splitterG8ton245n43_n245_8_( clk_6 , buf_splitterG8ton245n43_n245_7 , 0 , buf_splitterG8ton245n43_n245_8 );
buf_AQFP buf_splitterG8ton245n43_n245_9_( clk_8 , buf_splitterG8ton245n43_n245_8 , 0 , buf_splitterG8ton245n43_n245_9 );
buf_AQFP buf_splitterG8ton245n43_n245_10_( clk_2 , buf_splitterG8ton245n43_n245_9 , 0 , buf_splitterG8ton245n43_n245_10 );
buf_AQFP buf_splitterG8ton245n43_n245_11_( clk_3 , buf_splitterG8ton245n43_n245_10 , 0 , buf_splitterG8ton245n43_n245_11 );
buf_AQFP buf_splitterG8ton245n43_n245_12_( clk_5 , buf_splitterG8ton245n43_n245_11 , 0 , buf_splitterG8ton245n43_n245_12 );
buf_AQFP buf_splitterG8ton245n43_n246_1_( clk_8 , splitterG8ton245n43 , 0 , buf_splitterG8ton245n43_n246_1 );
buf_AQFP buf_splitterG8ton245n43_n246_2_( clk_2 , buf_splitterG8ton245n43_n246_1 , 0 , buf_splitterG8ton245n43_n246_2 );
buf_AQFP buf_splitterG8ton245n43_n246_3_( clk_4 , buf_splitterG8ton245n43_n246_2 , 0 , buf_splitterG8ton245n43_n246_3 );
buf_AQFP buf_splitterG8ton245n43_n246_4_( clk_6 , buf_splitterG8ton245n43_n246_3 , 0 , buf_splitterG8ton245n43_n246_4 );
buf_AQFP buf_splitterG8ton245n43_n246_5_( clk_8 , buf_splitterG8ton245n43_n246_4 , 0 , buf_splitterG8ton245n43_n246_5 );
buf_AQFP buf_splitterG8ton245n43_n246_6_( clk_2 , buf_splitterG8ton245n43_n246_5 , 0 , buf_splitterG8ton245n43_n246_6 );
buf_AQFP buf_splitterG8ton245n43_n246_7_( clk_4 , buf_splitterG8ton245n43_n246_6 , 0 , buf_splitterG8ton245n43_n246_7 );
buf_AQFP buf_splitterG8ton245n43_n246_8_( clk_6 , buf_splitterG8ton245n43_n246_7 , 0 , buf_splitterG8ton245n43_n246_8 );
buf_AQFP buf_splitterG8ton245n43_n246_9_( clk_8 , buf_splitterG8ton245n43_n246_8 , 0 , buf_splitterG8ton245n43_n246_9 );
buf_AQFP buf_splitterG8ton245n43_n246_10_( clk_2 , buf_splitterG8ton245n43_n246_9 , 0 , buf_splitterG8ton245n43_n246_10 );
buf_AQFP buf_splitterG8ton245n43_n246_11_( clk_4 , buf_splitterG8ton245n43_n246_10 , 0 , buf_splitterG8ton245n43_n246_11 );
buf_AQFP buf_splitterG8ton245n43_n246_12_( clk_6 , buf_splitterG8ton245n43_n246_11 , 0 , buf_splitterG8ton245n43_n246_12 );
buf_AQFP buf_splitterG9ton103n59_n249_1_( clk_5 , splitterG9ton103n59 , 0 , buf_splitterG9ton103n59_n249_1 );
buf_AQFP buf_splitterG9ton103n59_n249_2_( clk_7 , buf_splitterG9ton103n59_n249_1 , 0 , buf_splitterG9ton103n59_n249_2 );
buf_AQFP buf_splitterG9ton103n59_n249_3_( clk_1 , buf_splitterG9ton103n59_n249_2 , 0 , buf_splitterG9ton103n59_n249_3 );
buf_AQFP buf_splitterG9ton103n59_n249_4_( clk_3 , buf_splitterG9ton103n59_n249_3 , 0 , buf_splitterG9ton103n59_n249_4 );
buf_AQFP buf_splitterG9ton103n59_n249_5_( clk_5 , buf_splitterG9ton103n59_n249_4 , 0 , buf_splitterG9ton103n59_n249_5 );
buf_AQFP buf_splitterG9ton103n59_n249_6_( clk_7 , buf_splitterG9ton103n59_n249_5 , 0 , buf_splitterG9ton103n59_n249_6 );
buf_AQFP buf_splitterG9ton103n59_n249_7_( clk_1 , buf_splitterG9ton103n59_n249_6 , 0 , buf_splitterG9ton103n59_n249_7 );
buf_AQFP buf_splitterG9ton103n59_n249_8_( clk_3 , buf_splitterG9ton103n59_n249_7 , 0 , buf_splitterG9ton103n59_n249_8 );
buf_AQFP buf_splitterG9ton103n59_n249_9_( clk_5 , buf_splitterG9ton103n59_n249_8 , 0 , buf_splitterG9ton103n59_n249_9 );
buf_AQFP buf_splitterG9ton103n59_n249_10_( clk_7 , buf_splitterG9ton103n59_n249_9 , 0 , buf_splitterG9ton103n59_n249_10 );
buf_AQFP buf_splitterG9ton103n59_n249_11_( clk_1 , buf_splitterG9ton103n59_n249_10 , 0 , buf_splitterG9ton103n59_n249_11 );
buf_AQFP buf_splitterG9ton103n59_n249_12_( clk_3 , buf_splitterG9ton103n59_n249_11 , 0 , buf_splitterG9ton103n59_n249_12 );
buf_AQFP buf_splitterG9ton103n59_n249_13_( clk_5 , buf_splitterG9ton103n59_n249_12 , 0 , buf_splitterG9ton103n59_n249_13 );
buf_AQFP buf_splitterG9ton250n59_n250_1_( clk_2 , splitterG9ton250n59 , 0 , buf_splitterG9ton250n59_n250_1 );
buf_AQFP buf_splitterG9ton250n59_n250_2_( clk_4 , buf_splitterG9ton250n59_n250_1 , 0 , buf_splitterG9ton250n59_n250_2 );
buf_AQFP buf_splitterG9ton250n59_n250_3_( clk_6 , buf_splitterG9ton250n59_n250_2 , 0 , buf_splitterG9ton250n59_n250_3 );
buf_AQFP buf_splitterG9ton250n59_n250_4_( clk_7 , buf_splitterG9ton250n59_n250_3 , 0 , buf_splitterG9ton250n59_n250_4 );
buf_AQFP buf_splitterG9ton250n59_n250_5_( clk_8 , buf_splitterG9ton250n59_n250_4 , 0 , buf_splitterG9ton250n59_n250_5 );
buf_AQFP buf_splitterG9ton250n59_n250_6_( clk_2 , buf_splitterG9ton250n59_n250_5 , 0 , buf_splitterG9ton250n59_n250_6 );
buf_AQFP buf_splitterG9ton250n59_n250_7_( clk_4 , buf_splitterG9ton250n59_n250_6 , 0 , buf_splitterG9ton250n59_n250_7 );
buf_AQFP buf_splitterG9ton250n59_n250_8_( clk_6 , buf_splitterG9ton250n59_n250_7 , 0 , buf_splitterG9ton250n59_n250_8 );
buf_AQFP buf_splitterG9ton250n59_n250_9_( clk_8 , buf_splitterG9ton250n59_n250_8 , 0 , buf_splitterG9ton250n59_n250_9 );
buf_AQFP buf_splitterG9ton250n59_n250_10_( clk_2 , buf_splitterG9ton250n59_n250_9 , 0 , buf_splitterG9ton250n59_n250_10 );
buf_AQFP buf_splitterG9ton250n59_n250_11_( clk_4 , buf_splitterG9ton250n59_n250_10 , 0 , buf_splitterG9ton250n59_n250_11 );
buf_AQFP buf_splitterfromn34_n74_1_( clk_6 , splitterfromn34 , 0 , buf_splitterfromn34_n74_1 );
buf_AQFP buf_splittern35ton252n78_n252_1_( clk_6 , splittern35ton252n78 , 0 , buf_splittern35ton252n78_n252_1 );
buf_AQFP buf_splittern35ton252n78_n252_2_( clk_8 , buf_splittern35ton252n78_n252_1 , 0 , buf_splittern35ton252n78_n252_2 );
buf_AQFP buf_splittern35ton252n78_n78_1_( clk_6 , splittern35ton252n78 , 0 , buf_splittern35ton252n78_n78_1 );
buf_AQFP buf_splittern41ton54n94_n54_1_( clk_4 , splittern41ton54n94 , 0 , buf_splittern41ton54n94_n54_1 );
buf_AQFP buf_splittern41ton54n94_n55_1_( clk_4 , splittern41ton54n94 , 0 , buf_splittern41ton54n94_n55_1 );
buf_AQFP buf_splittern50ton186n52_n186_1_( clk_2 , splittern50ton186n52 , 0 , buf_splittern50ton186n52_n186_1 );
buf_AQFP buf_splittern50ton186n52_n187_1_( clk_2 , splittern50ton186n52 , 0 , buf_splittern50ton186n52_n187_1 );
buf_AQFP buf_splittern66ton67n86_n67_1_( clk_3 , splittern66ton67n86 , 0 , buf_splittern66ton67n86_n67_1 );
buf_AQFP buf_splittern66ton67n86_n68_1_( clk_3 , splittern66ton67n86 , 0 , buf_splittern66ton67n86_n68_1 );
buf_AQFP buf_splitterfromn72_n277_1_( clk_4 , splitterfromn72 , 0 , buf_splitterfromn72_n277_1 );
buf_AQFP buf_splitterfromn72_n277_2_( clk_6 , buf_splitterfromn72_n277_1 , 0 , buf_splitterfromn72_n277_2 );
buf_AQFP buf_splitterfromn72_n277_3_( clk_8 , buf_splitterfromn72_n277_2 , 0 , buf_splitterfromn72_n277_3 );
buf_AQFP buf_splitterfromn72_n277_4_( clk_2 , buf_splitterfromn72_n277_3 , 0 , buf_splitterfromn72_n277_4 );
buf_AQFP buf_splitterfromn72_n277_5_( clk_4 , buf_splitterfromn72_n277_4 , 0 , buf_splitterfromn72_n277_5 );
buf_AQFP buf_splitterfromn72_n277_6_( clk_6 , buf_splitterfromn72_n277_5 , 0 , buf_splitterfromn72_n277_6 );
buf_AQFP buf_splitterfromn72_n277_7_( clk_8 , buf_splitterfromn72_n277_6 , 0 , buf_splitterfromn72_n277_7 );
buf_AQFP buf_splitterfromn72_n277_8_( clk_1 , buf_splitterfromn72_n277_7 , 0 , buf_splitterfromn72_n277_8 );
buf_AQFP buf_splitterfromn72_n277_9_( clk_3 , buf_splitterfromn72_n277_8 , 0 , buf_splitterfromn72_n277_9 );
buf_AQFP buf_splittern73ton278n76_n278_1_( clk_5 , splittern73ton278n76 , 0 , buf_splittern73ton278n76_n278_1 );
buf_AQFP buf_splittern73ton278n76_n278_2_( clk_7 , buf_splittern73ton278n76_n278_1 , 0 , buf_splittern73ton278n76_n278_2 );
buf_AQFP buf_splittern73ton278n76_n278_3_( clk_1 , buf_splittern73ton278n76_n278_2 , 0 , buf_splittern73ton278n76_n278_3 );
buf_AQFP buf_splittern73ton278n76_n278_4_( clk_3 , buf_splittern73ton278n76_n278_3 , 0 , buf_splittern73ton278n76_n278_4 );
buf_AQFP buf_splittern73ton278n76_n278_5_( clk_5 , buf_splittern73ton278n76_n278_4 , 0 , buf_splittern73ton278n76_n278_5 );
buf_AQFP buf_splittern73ton278n76_n278_6_( clk_7 , buf_splittern73ton278n76_n278_5 , 0 , buf_splittern73ton278n76_n278_6 );
buf_AQFP buf_splittern73ton278n76_n278_7_( clk_1 , buf_splittern73ton278n76_n278_6 , 0 , buf_splittern73ton278n76_n278_7 );
buf_AQFP buf_splittern74ton275n76_n275_1_( clk_4 , splittern74ton275n76 , 0 , buf_splittern74ton275n76_n275_1 );
buf_AQFP buf_splittern74ton275n76_n275_2_( clk_5 , buf_splittern74ton275n76_n275_1 , 0 , buf_splittern74ton275n76_n275_2 );
buf_AQFP buf_splittern74ton275n76_n275_3_( clk_7 , buf_splittern74ton275n76_n275_2 , 0 , buf_splittern74ton275n76_n275_3 );
buf_AQFP buf_splittern74ton275n76_n275_4_( clk_1 , buf_splittern74ton275n76_n275_3 , 0 , buf_splittern74ton275n76_n275_4 );
buf_AQFP buf_splittern74ton275n76_n275_5_( clk_3 , buf_splittern74ton275n76_n275_4 , 0 , buf_splittern74ton275n76_n275_5 );
buf_AQFP buf_splittern74ton275n76_n275_6_( clk_4 , buf_splittern74ton275n76_n275_5 , 0 , buf_splittern74ton275n76_n275_6 );
buf_AQFP buf_splittern74ton275n76_n275_7_( clk_6 , buf_splittern74ton275n76_n275_6 , 0 , buf_splittern74ton275n76_n275_7 );
buf_AQFP buf_splittern74ton275n76_n275_8_( clk_8 , buf_splittern74ton275n76_n275_7 , 0 , buf_splittern74ton275n76_n275_8 );
buf_AQFP buf_splittern77ton253n78_n253_1_( clk_1 , splittern77ton253n78 , 0 , buf_splittern77ton253n78_n253_1 );
buf_AQFP buf_splittern87ton189n97_n189_1_( clk_6 , splittern87ton189n97 , 0 , buf_splittern87ton189n97_n189_1 );
buf_AQFP buf_splittern87ton189n97_n190_1_( clk_5 , splittern87ton189n97 , 0 , buf_splittern87ton189n97_n190_1 );
buf_AQFP buf_splitterfromn98_n321_1_( clk_1 , splitterfromn98 , 0 , buf_splitterfromn98_n321_1 );
buf_AQFP buf_splitterfromn98_n321_2_( clk_2 , buf_splitterfromn98_n321_1 , 0 , buf_splitterfromn98_n321_2 );
buf_AQFP buf_splitterfromn98_n321_3_( clk_3 , buf_splitterfromn98_n321_2 , 0 , buf_splitterfromn98_n321_3 );
buf_AQFP buf_splitterfromn98_n321_4_( clk_5 , buf_splitterfromn98_n321_3 , 0 , buf_splitterfromn98_n321_4 );
buf_AQFP buf_splitterfromn98_n321_5_( clk_7 , buf_splitterfromn98_n321_4 , 0 , buf_splitterfromn98_n321_5 );
buf_AQFP buf_splitterfromn98_n321_6_( clk_1 , buf_splitterfromn98_n321_5 , 0 , buf_splitterfromn98_n321_6 );
buf_AQFP buf_splitterfromn98_n321_7_( clk_3 , buf_splitterfromn98_n321_6 , 0 , buf_splitterfromn98_n321_7 );
buf_AQFP buf_splitterfromn98_n321_8_( clk_5 , buf_splitterfromn98_n321_7 , 0 , buf_splitterfromn98_n321_8 );
buf_AQFP buf_splitterfromn98_n321_9_( clk_7 , buf_splitterfromn98_n321_8 , 0 , buf_splitterfromn98_n321_9 );
buf_AQFP buf_splitterfromn98_n321_10_( clk_1 , buf_splitterfromn98_n321_9 , 0 , buf_splitterfromn98_n321_10 );
buf_AQFP buf_splittern105ton106n309_n308_1_( clk_8 , splittern105ton106n309 , 0 , buf_splittern105ton106n309_n308_1 );
buf_AQFP buf_splittern105ton106n309_n308_2_( clk_1 , buf_splittern105ton106n309_n308_1 , 0 , buf_splittern105ton106n309_n308_2 );
buf_AQFP buf_splittern105ton106n309_n308_3_( clk_3 , buf_splittern105ton106n309_n308_2 , 0 , buf_splittern105ton106n309_n308_3 );
buf_AQFP buf_splittern105ton106n309_n309_1_( clk_8 , splittern105ton106n309 , 0 , buf_splittern105ton106n309_n309_1 );
buf_AQFP buf_splittern105ton106n309_n309_2_( clk_2 , buf_splittern105ton106n309_n309_1 , 0 , buf_splittern105ton106n309_n309_2 );
buf_AQFP buf_splittern105ton106n309_n309_3_( clk_3 , buf_splittern105ton106n309_n309_2 , 0 , buf_splittern105ton106n309_n309_3 );
buf_AQFP buf_splittern105ton106n309_n309_4_( clk_5 , buf_splittern105ton106n309_n309_3 , 0 , buf_splittern105ton106n309_n309_4 );
buf_AQFP buf_splitterfromn125_n297_1_( clk_2 , splitterfromn125 , 0 , buf_splitterfromn125_n297_1 );
buf_AQFP buf_splitterfromn125_n297_2_( clk_4 , buf_splitterfromn125_n297_1 , 0 , buf_splitterfromn125_n297_2 );
buf_AQFP buf_splitterfromn125_n297_3_( clk_6 , buf_splitterfromn125_n297_2 , 0 , buf_splitterfromn125_n297_3 );
buf_AQFP buf_splitterfromn125_n297_4_( clk_8 , buf_splitterfromn125_n297_3 , 0 , buf_splitterfromn125_n297_4 );
buf_AQFP buf_splitterfromn125_n297_5_( clk_2 , buf_splitterfromn125_n297_4 , 0 , buf_splitterfromn125_n297_5 );
buf_AQFP buf_splitterfromn125_n297_6_( clk_4 , buf_splitterfromn125_n297_5 , 0 , buf_splitterfromn125_n297_6 );
buf_AQFP buf_splitterfromn125_n297_7_( clk_5 , buf_splitterfromn125_n297_6 , 0 , buf_splitterfromn125_n297_7 );
buf_AQFP buf_splitterfromn125_n297_8_( clk_6 , buf_splitterfromn125_n297_7 , 0 , buf_splitterfromn125_n297_8 );
buf_AQFP buf_splitterfromn125_n297_9_( clk_8 , buf_splitterfromn125_n297_8 , 0 , buf_splitterfromn125_n297_9 );
buf_AQFP buf_splitterfromn125_n297_10_( clk_1 , buf_splitterfromn125_n297_9 , 0 , buf_splitterfromn125_n297_10 );
buf_AQFP buf_splittern128ton129n295_n295_1_( clk_4 , splittern128ton129n295 , 0 , buf_splittern128ton129n295_n295_1 );
buf_AQFP buf_splitterfromn151_n289_1_( clk_2 , splitterfromn151 , 0 , buf_splitterfromn151_n289_1 );
buf_AQFP buf_splitterfromn151_n289_2_( clk_4 , buf_splitterfromn151_n289_1 , 0 , buf_splitterfromn151_n289_2 );
buf_AQFP buf_splitterfromn151_n289_3_( clk_6 , buf_splitterfromn151_n289_2 , 0 , buf_splitterfromn151_n289_3 );
buf_AQFP buf_splitterfromn151_n289_4_( clk_8 , buf_splitterfromn151_n289_3 , 0 , buf_splitterfromn151_n289_4 );
buf_AQFP buf_splitterfromn151_n289_5_( clk_2 , buf_splitterfromn151_n289_4 , 0 , buf_splitterfromn151_n289_5 );
buf_AQFP buf_splitterfromn151_n289_6_( clk_4 , buf_splitterfromn151_n289_5 , 0 , buf_splitterfromn151_n289_6 );
buf_AQFP buf_splitterfromn151_n289_7_( clk_6 , buf_splitterfromn151_n289_6 , 0 , buf_splitterfromn151_n289_7 );
buf_AQFP buf_splitterfromn151_n289_8_( clk_8 , buf_splitterfromn151_n289_7 , 0 , buf_splitterfromn151_n289_8 );
buf_AQFP buf_splitterfromn151_n289_9_( clk_2 , buf_splitterfromn151_n289_8 , 0 , buf_splitterfromn151_n289_9 );
buf_AQFP buf_splitterfromn171_n293_1_( clk_2 , splitterfromn171 , 0 , buf_splitterfromn171_n293_1 );
buf_AQFP buf_splitterfromn171_n293_2_( clk_4 , buf_splitterfromn171_n293_1 , 0 , buf_splitterfromn171_n293_2 );
buf_AQFP buf_splitterfromn171_n293_3_( clk_6 , buf_splitterfromn171_n293_2 , 0 , buf_splitterfromn171_n293_3 );
buf_AQFP buf_splitterfromn171_n293_4_( clk_8 , buf_splitterfromn171_n293_3 , 0 , buf_splitterfromn171_n293_4 );
buf_AQFP buf_splitterfromn171_n293_5_( clk_2 , buf_splitterfromn171_n293_4 , 0 , buf_splitterfromn171_n293_5 );
buf_AQFP buf_splitterfromn171_n293_6_( clk_4 , buf_splitterfromn171_n293_5 , 0 , buf_splitterfromn171_n293_6 );
buf_AQFP buf_splitterfromn171_n293_7_( clk_6 , buf_splitterfromn171_n293_6 , 0 , buf_splitterfromn171_n293_7 );
buf_AQFP buf_splitterfromn171_n293_8_( clk_8 , buf_splitterfromn171_n293_7 , 0 , buf_splitterfromn171_n293_8 );
buf_AQFP buf_splitterfromn171_n293_9_( clk_2 , buf_splitterfromn171_n293_8 , 0 , buf_splitterfromn171_n293_9 );
buf_AQFP buf_splittern177ton197n272_n272_1_( clk_8 , splittern177ton197n272 , 0 , buf_splittern177ton197n272_n272_1 );
buf_AQFP buf_splitterfromn191_n283_1_( clk_2 , splitterfromn191 , 0 , buf_splitterfromn191_n283_1 );
buf_AQFP buf_splitterfromn191_n283_2_( clk_3 , buf_splitterfromn191_n283_1 , 0 , buf_splitterfromn191_n283_2 );
buf_AQFP buf_splitterfromn191_n283_3_( clk_5 , buf_splitterfromn191_n283_2 , 0 , buf_splitterfromn191_n283_3 );
buf_AQFP buf_splitterfromn191_n283_4_( clk_7 , buf_splitterfromn191_n283_3 , 0 , buf_splitterfromn191_n283_4 );
buf_AQFP buf_splitterfromn191_n283_5_( clk_1 , buf_splitterfromn191_n283_4 , 0 , buf_splitterfromn191_n283_5 );
buf_AQFP buf_splitterfromn191_n283_6_( clk_3 , buf_splitterfromn191_n283_5 , 0 , buf_splitterfromn191_n283_6 );
buf_AQFP buf_splitterfromn191_n283_7_( clk_5 , buf_splitterfromn191_n283_6 , 0 , buf_splitterfromn191_n283_7 );
buf_AQFP buf_splitterfromn191_n283_8_( clk_7 , buf_splitterfromn191_n283_7 , 0 , buf_splitterfromn191_n283_8 );
buf_AQFP buf_splitterfromn191_n283_9_( clk_1 , buf_splitterfromn191_n283_8 , 0 , buf_splitterfromn191_n283_9 );
buf_AQFP buf_splitterfromn191_n283_10_( clk_3 , buf_splitterfromn191_n283_9 , 0 , buf_splitterfromn191_n283_10 );
buf_AQFP buf_splittern192ton193n284_n284_1_( clk_5 , splittern192ton193n284 , 0 , buf_splittern192ton193n284_n284_1 );
buf_AQFP buf_splittern192ton193n284_n284_2_( clk_7 , buf_splittern192ton193n284_n284_1 , 0 , buf_splittern192ton193n284_n284_2 );
buf_AQFP buf_splittern192ton193n284_n284_3_( clk_1 , buf_splittern192ton193n284_n284_2 , 0 , buf_splittern192ton193n284_n284_3 );
buf_AQFP buf_splittern192ton193n284_n284_4_( clk_3 , buf_splittern192ton193n284_n284_3 , 0 , buf_splittern192ton193n284_n284_4 );
buf_AQFP buf_splittern192ton193n284_n284_5_( clk_5 , buf_splittern192ton193n284_n284_4 , 0 , buf_splittern192ton193n284_n284_5 );
buf_AQFP buf_splittern192ton193n284_n284_6_( clk_7 , buf_splittern192ton193n284_n284_5 , 0 , buf_splittern192ton193n284_n284_6 );
buf_AQFP buf_splittern192ton193n284_n284_7_( clk_1 , buf_splittern192ton193n284_n284_6 , 0 , buf_splittern192ton193n284_n284_7 );
buf_AQFP buf_splitterfromn200_n204_1_( clk_6 , splitterfromn200 , 0 , buf_splitterfromn200_n204_1 );
buf_AQFP buf_splittern203ton204n321_n279_1_( clk_8 , splittern203ton204n321 , 0 , buf_splittern203ton204n321_n279_1 );
buf_AQFP buf_splittern203ton204n321_n279_2_( clk_2 , buf_splittern203ton204n321_n279_1 , 0 , buf_splittern203ton204n321_n279_2 );
buf_AQFP buf_splittern203ton204n321_n279_3_( clk_4 , buf_splittern203ton204n321_n279_2 , 0 , buf_splittern203ton204n321_n279_3 );
buf_AQFP buf_splittern203ton204n321_n279_4_( clk_6 , buf_splittern203ton204n321_n279_3 , 0 , buf_splittern203ton204n321_n279_4 );
buf_AQFP buf_splittern203ton204n321_n279_5_( clk_7 , buf_splittern203ton204n321_n279_4 , 0 , buf_splittern203ton204n321_n279_5 );
buf_AQFP buf_splittern203ton204n321_n279_6_( clk_8 , buf_splittern203ton204n321_n279_5 , 0 , buf_splittern203ton204n321_n279_6 );
buf_AQFP buf_splittern203ton204n321_n279_7_( clk_1 , buf_splittern203ton204n321_n279_6 , 0 , buf_splittern203ton204n321_n279_7 );
buf_AQFP buf_splittern203ton204n321_n279_8_( clk_2 , buf_splittern203ton204n321_n279_7 , 0 , buf_splittern203ton204n321_n279_8 );
buf_AQFP buf_splittern203ton204n321_n279_9_( clk_4 , buf_splittern203ton204n321_n279_8 , 0 , buf_splittern203ton204n321_n279_9 );
buf_AQFP buf_splittern203ton204n321_n279_10_( clk_5 , buf_splittern203ton204n321_n279_9 , 0 , buf_splittern203ton204n321_n279_10 );
buf_AQFP buf_splittern203ton204n321_n279_11_( clk_7 , buf_splittern203ton204n321_n279_10 , 0 , buf_splittern203ton204n321_n279_11 );
buf_AQFP buf_splittern203ton204n321_n279_12_( clk_1 , buf_splittern203ton204n321_n279_11 , 0 , buf_splittern203ton204n321_n279_12 );
buf_AQFP buf_splittern203ton204n321_n279_13_( clk_3 , buf_splittern203ton204n321_n279_12 , 0 , buf_splittern203ton204n321_n279_13 );
buf_AQFP buf_splittern203ton204n321_n285_1_( clk_8 , splittern203ton204n321 , 0 , buf_splittern203ton204n321_n285_1 );
buf_AQFP buf_splittern203ton204n321_n285_2_( clk_2 , buf_splittern203ton204n321_n285_1 , 0 , buf_splittern203ton204n321_n285_2 );
buf_AQFP buf_splittern203ton204n321_n285_3_( clk_3 , buf_splittern203ton204n321_n285_2 , 0 , buf_splittern203ton204n321_n285_3 );
buf_AQFP buf_splittern203ton204n321_n285_4_( clk_4 , buf_splittern203ton204n321_n285_3 , 0 , buf_splittern203ton204n321_n285_4 );
buf_AQFP buf_splittern203ton204n321_n285_5_( clk_5 , buf_splittern203ton204n321_n285_4 , 0 , buf_splittern203ton204n321_n285_5 );
buf_AQFP buf_splittern203ton204n321_n285_6_( clk_7 , buf_splittern203ton204n321_n285_5 , 0 , buf_splittern203ton204n321_n285_6 );
buf_AQFP buf_splittern203ton204n321_n285_7_( clk_8 , buf_splittern203ton204n321_n285_6 , 0 , buf_splittern203ton204n321_n285_7 );
buf_AQFP buf_splittern203ton204n321_n285_8_( clk_2 , buf_splittern203ton204n321_n285_7 , 0 , buf_splittern203ton204n321_n285_8 );
buf_AQFP buf_splittern203ton204n321_n285_9_( clk_3 , buf_splittern203ton204n321_n285_8 , 0 , buf_splittern203ton204n321_n285_9 );
buf_AQFP buf_splittern203ton204n321_n285_10_( clk_4 , buf_splittern203ton204n321_n285_9 , 0 , buf_splittern203ton204n321_n285_10 );
buf_AQFP buf_splittern203ton204n321_n285_11_( clk_5 , buf_splittern203ton204n321_n285_10 , 0 , buf_splittern203ton204n321_n285_11 );
buf_AQFP buf_splittern203ton204n321_n285_12_( clk_7 , buf_splittern203ton204n321_n285_11 , 0 , buf_splittern203ton204n321_n285_12 );
buf_AQFP buf_splittern203ton204n321_n285_13_( clk_1 , buf_splittern203ton204n321_n285_12 , 0 , buf_splittern203ton204n321_n285_13 );
buf_AQFP buf_splittern203ton204n321_n285_14_( clk_3 , buf_splittern203ton204n321_n285_13 , 0 , buf_splittern203ton204n321_n285_14 );
buf_AQFP buf_splittern203ton290n321_n290_1_( clk_3 , splittern203ton290n321 , 0 , buf_splittern203ton290n321_n290_1 );
buf_AQFP buf_splittern203ton290n321_n294_1_( clk_3 , splittern203ton290n321 , 0 , buf_splittern203ton290n321_n294_1 );
buf_AQFP buf_splitterfromn205_n206_1_( clk_5 , splitterfromn205 , 0 , buf_splitterfromn205_n206_1 );
buf_AQFP buf_splitterfromn205_n206_2_( clk_7 , buf_splitterfromn205_n206_1 , 0 , buf_splitterfromn205_n206_2 );
buf_AQFP buf_splitterfromn205_n206_3_( clk_8 , buf_splitterfromn205_n206_2 , 0 , buf_splitterfromn205_n206_3 );
buf_AQFP buf_splitterfromn205_n206_4_( clk_2 , buf_splitterfromn205_n206_3 , 0 , buf_splitterfromn205_n206_4 );
buf_AQFP buf_splitterfromn205_n235_1_( clk_5 , splitterfromn205 , 0 , buf_splitterfromn205_n235_1 );
buf_AQFP buf_splitterfromn205_n235_2_( clk_6 , buf_splitterfromn205_n235_1 , 0 , buf_splitterfromn205_n235_2 );
buf_AQFP buf_splitterfromn205_n235_3_( clk_7 , buf_splitterfromn205_n235_2 , 0 , buf_splitterfromn205_n235_3 );
buf_AQFP buf_splitterfromn205_n235_4_( clk_8 , buf_splitterfromn205_n235_3 , 0 , buf_splitterfromn205_n235_4 );
buf_AQFP buf_splitterfromn205_n235_5_( clk_1 , buf_splitterfromn205_n235_4 , 0 , buf_splitterfromn205_n235_5 );
buf_AQFP buf_splitterfromn205_n235_6_( clk_2 , buf_splitterfromn205_n235_5 , 0 , buf_splitterfromn205_n235_6 );
buf_AQFP buf_splitterfromn219_n310_1_( clk_8 , splitterfromn219 , 0 , buf_splitterfromn219_n310_1 );
buf_AQFP buf_splittern221ton222n254_n222_1_( clk_1 , splittern221ton222n254 , 0 , buf_splittern221ton222n254_n222_1 );
buf_AQFP buf_splittern221ton222n254_n222_2_( clk_3 , buf_splittern221ton222n254_n222_1 , 0 , buf_splittern221ton222n254_n222_2 );
buf_AQFP buf_splittern221ton222n254_n248_1_( clk_1 , splittern221ton222n254 , 0 , buf_splittern221ton222n254_n248_1 );
buf_AQFP buf_splittern221ton222n254_n248_2_( clk_2 , buf_splittern221ton222n254_n248_1 , 0 , buf_splittern221ton222n254_n248_2 );
buf_AQFP buf_splittern221ton222n254_n254_1_( clk_1 , splittern221ton222n254 , 0 , buf_splittern221ton222n254_n254_1 );
buf_AQFP buf_splittern221ton222n254_n254_2_( clk_3 , buf_splittern221ton222n254_n254_1 , 0 , buf_splittern221ton222n254_n254_2 );
buf_AQFP buf_splitterfromn299_n305_1_( clk_3 , splitterfromn299 , 0 , buf_splitterfromn299_n305_1 );
buf_AQFP buf_splitterfromn299_n305_2_( clk_5 , buf_splitterfromn299_n305_1 , 0 , buf_splitterfromn299_n305_2 );
buf_AQFP buf_splitterfromn299_n305_3_( clk_7 , buf_splitterfromn299_n305_2 , 0 , buf_splitterfromn299_n305_3 );
buf_AQFP buf_splitterfromn299_n305_4_( clk_1 , buf_splitterfromn299_n305_3 , 0 , buf_splitterfromn299_n305_4 );
buf_AQFP buf_splitterfromn299_n305_5_( clk_3 , buf_splitterfromn299_n305_4 , 0 , buf_splitterfromn299_n305_5 );
buf_AQFP buf_splitterfromn299_n305_6_( clk_5 , buf_splitterfromn299_n305_5 , 0 , buf_splitterfromn299_n305_6 );
buf_AQFP buf_splitterfromn299_n305_7_( clk_7 , buf_splitterfromn299_n305_6 , 0 , buf_splitterfromn299_n305_7 );
buf_AQFP buf_splitterfromn299_n305_8_( clk_1 , buf_splitterfromn299_n305_7 , 0 , buf_splitterfromn299_n305_8 );
buf_AQFP buf_splitterfromn299_n306_1_( clk_3 , splitterfromn299 , 0 , buf_splitterfromn299_n306_1 );
buf_AQFP buf_splitterfromn299_n306_2_( clk_5 , buf_splitterfromn299_n306_1 , 0 , buf_splitterfromn299_n306_2 );
buf_AQFP buf_splitterfromn299_n306_3_( clk_7 , buf_splitterfromn299_n306_2 , 0 , buf_splitterfromn299_n306_3 );
buf_AQFP buf_splitterfromn299_n306_4_( clk_1 , buf_splitterfromn299_n306_3 , 0 , buf_splitterfromn299_n306_4 );
buf_AQFP buf_splitterfromn299_n306_5_( clk_3 , buf_splitterfromn299_n306_4 , 0 , buf_splitterfromn299_n306_5 );
buf_AQFP buf_splitterfromn299_n306_6_( clk_5 , buf_splitterfromn299_n306_5 , 0 , buf_splitterfromn299_n306_6 );
buf_AQFP buf_splitterfromn299_n306_7_( clk_7 , buf_splitterfromn299_n306_6 , 0 , buf_splitterfromn299_n306_7 );
buf_AQFP buf_splitterfromn299_n306_8_( clk_1 , buf_splitterfromn299_n306_7 , 0 , buf_splitterfromn299_n306_8 );
buf_AQFP buf_splitterfromn300_n301_1_( clk_8 , splitterfromn300 , 0 , buf_splitterfromn300_n301_1 );
buf_AQFP buf_splitterfromn300_n301_2_( clk_2 , buf_splitterfromn300_n301_1 , 0 , buf_splitterfromn300_n301_2 );
buf_AQFP buf_splitterfromn300_n301_3_( clk_4 , buf_splitterfromn300_n301_2 , 0 , buf_splitterfromn300_n301_3 );
buf_AQFP buf_splitterfromn300_n301_4_( clk_6 , buf_splitterfromn300_n301_3 , 0 , buf_splitterfromn300_n301_4 );
buf_AQFP buf_splitterfromn300_n301_5_( clk_7 , buf_splitterfromn300_n301_4 , 0 , buf_splitterfromn300_n301_5 );
buf_AQFP buf_splitterfromn300_n301_6_( clk_8 , buf_splitterfromn300_n301_5 , 0 , buf_splitterfromn300_n301_6 );
buf_AQFP buf_splitterfromn300_n301_7_( clk_2 , buf_splitterfromn300_n301_6 , 0 , buf_splitterfromn300_n301_7 );
buf_AQFP buf_splitterfromn300_n301_8_( clk_3 , buf_splitterfromn300_n301_7 , 0 , buf_splitterfromn300_n301_8 );
buf_AQFP buf_splitterfromn300_n301_9_( clk_5 , buf_splitterfromn300_n301_8 , 0 , buf_splitterfromn300_n301_9 );
buf_AQFP buf_splitterfromn300_n302_1_( clk_7 , splitterfromn300 , 0 , buf_splitterfromn300_n302_1 );
buf_AQFP buf_splitterfromn300_n302_2_( clk_8 , buf_splitterfromn300_n302_1 , 0 , buf_splitterfromn300_n302_2 );
buf_AQFP buf_splitterfromn300_n302_3_( clk_1 , buf_splitterfromn300_n302_2 , 0 , buf_splitterfromn300_n302_3 );
buf_AQFP buf_splitterfromn300_n302_4_( clk_3 , buf_splitterfromn300_n302_3 , 0 , buf_splitterfromn300_n302_4 );
buf_AQFP buf_splitterfromn300_n302_5_( clk_4 , buf_splitterfromn300_n302_4 , 0 , buf_splitterfromn300_n302_5 );
buf_AQFP buf_splitterfromn300_n302_6_( clk_5 , buf_splitterfromn300_n302_5 , 0 , buf_splitterfromn300_n302_6 );
buf_AQFP buf_splitterfromn300_n302_7_( clk_7 , buf_splitterfromn300_n302_6 , 0 , buf_splitterfromn300_n302_7 );
buf_AQFP buf_splitterfromn300_n302_8_( clk_1 , buf_splitterfromn300_n302_7 , 0 , buf_splitterfromn300_n302_8 );
buf_AQFP buf_splitterfromn300_n302_9_( clk_3 , buf_splitterfromn300_n302_8 , 0 , buf_splitterfromn300_n302_9 );
buf_AQFP buf_splitterfromn300_n302_10_( clk_5 , buf_splitterfromn300_n302_9 , 0 , buf_splitterfromn300_n302_10 );
buf_AQFP buf_splitterfromn311_n317_1_( clk_5 , splitterfromn311 , 0 , buf_splitterfromn311_n317_1 );
buf_AQFP buf_splitterfromn311_n317_2_( clk_7 , buf_splitterfromn311_n317_1 , 0 , buf_splitterfromn311_n317_2 );
buf_AQFP buf_splitterfromn311_n317_3_( clk_1 , buf_splitterfromn311_n317_2 , 0 , buf_splitterfromn311_n317_3 );
buf_AQFP buf_splitterfromn311_n318_1_( clk_4 , splitterfromn311 , 0 , buf_splitterfromn311_n318_1 );
buf_AQFP buf_splitterfromn311_n318_2_( clk_5 , buf_splitterfromn311_n318_1 , 0 , buf_splitterfromn311_n318_2 );
buf_AQFP buf_splitterfromn311_n318_3_( clk_7 , buf_splitterfromn311_n318_2 , 0 , buf_splitterfromn311_n318_3 );
buf_AQFP buf_splitterfromn311_n318_4_( clk_1 , buf_splitterfromn311_n318_3 , 0 , buf_splitterfromn311_n318_4 );
buf_AQFP buf_splitterfromn312_n313_1_( clk_7 , splitterfromn312 , 0 , buf_splitterfromn312_n313_1 );
buf_AQFP buf_splitterfromn312_n313_2_( clk_8 , buf_splitterfromn312_n313_1 , 0 , buf_splitterfromn312_n313_2 );
buf_AQFP buf_splitterfromn312_n313_3_( clk_2 , buf_splitterfromn312_n313_2 , 0 , buf_splitterfromn312_n313_3 );
buf_AQFP buf_splitterfromn312_n313_4_( clk_4 , buf_splitterfromn312_n313_3 , 0 , buf_splitterfromn312_n313_4 );
buf_AQFP buf_splitterfromn312_n313_5_( clk_6 , buf_splitterfromn312_n313_4 , 0 , buf_splitterfromn312_n313_5 );
buf_AQFP buf_splitterfromn312_n313_6_( clk_7 , buf_splitterfromn312_n313_5 , 0 , buf_splitterfromn312_n313_6 );
buf_AQFP buf_splitterfromn312_n313_7_( clk_1 , buf_splitterfromn312_n313_6 , 0 , buf_splitterfromn312_n313_7 );
buf_AQFP buf_splitterfromn312_n313_8_( clk_2 , buf_splitterfromn312_n313_7 , 0 , buf_splitterfromn312_n313_8 );
buf_AQFP buf_splitterfromn312_n313_9_( clk_3 , buf_splitterfromn312_n313_8 , 0 , buf_splitterfromn312_n313_9 );
buf_AQFP buf_splitterfromn312_n313_10_( clk_5 , buf_splitterfromn312_n313_9 , 0 , buf_splitterfromn312_n313_10 );
buf_AQFP buf_splitterfromn312_n314_1_( clk_7 , splitterfromn312 , 0 , buf_splitterfromn312_n314_1 );
buf_AQFP buf_splitterfromn312_n314_2_( clk_8 , buf_splitterfromn312_n314_1 , 0 , buf_splitterfromn312_n314_2 );
buf_AQFP buf_splitterfromn312_n314_3_( clk_1 , buf_splitterfromn312_n314_2 , 0 , buf_splitterfromn312_n314_3 );
buf_AQFP buf_splitterfromn312_n314_4_( clk_2 , buf_splitterfromn312_n314_3 , 0 , buf_splitterfromn312_n314_4 );
buf_AQFP buf_splitterfromn312_n314_5_( clk_3 , buf_splitterfromn312_n314_4 , 0 , buf_splitterfromn312_n314_5 );
buf_AQFP buf_splitterfromn312_n314_6_( clk_4 , buf_splitterfromn312_n314_5 , 0 , buf_splitterfromn312_n314_6 );
buf_AQFP buf_splitterfromn312_n314_7_( clk_5 , buf_splitterfromn312_n314_6 , 0 , buf_splitterfromn312_n314_7 );
buf_AQFP buf_splitterfromn312_n314_8_( clk_6 , buf_splitterfromn312_n314_7 , 0 , buf_splitterfromn312_n314_8 );
buf_AQFP buf_splitterfromn312_n314_9_( clk_8 , buf_splitterfromn312_n314_8 , 0 , buf_splitterfromn312_n314_9 );
buf_AQFP buf_splitterfromn312_n314_10_( clk_2 , buf_splitterfromn312_n314_9 , 0 , buf_splitterfromn312_n314_10 );
buf_AQFP buf_splitterfromn312_n314_11_( clk_4 , buf_splitterfromn312_n314_10 , 0 , buf_splitterfromn312_n314_11 );
buf_AQFP buf_splitterfromn312_n314_12_( clk_5 , buf_splitterfromn312_n314_11 , 0 , buf_splitterfromn312_n314_12 );
splitter_AQFP splitterG1ton207n91_( clk_5 , buf_G1_splitterG1ton207n91_2 , 0 , splitterG1ton207n91 );
splitter_AQFP splitterG1ton49n91_( clk_6 , splitterG1ton207n91 , 0 , splitterG1ton49n91 );
splitter_AQFP splitterG10ton120n62_( clk_2 , G10 , 0 , splitterG10ton120n62 );
splitter_AQFP splitterG10ton224n62_( clk_3 , splitterG10ton120n62 , 0 , splitterG10ton224n62 );
splitter_AQFP splitterG11ton134n80_( clk_2 , G11 , 0 , splitterG11ton134n80 );
splitter_AQFP splitterG11ton256n80_( clk_3 , splitterG11ton134n80 , 0 , splitterG11ton256n80 );
splitter_AQFP splitterG12ton163n83_( clk_5 , buf_G12_splitterG12ton163n83_1 , 0 , splitterG12ton163n83 );
splitter_AQFP splitterG12ton259n83_( clk_6 , splitterG12ton163n83 , 0 , splitterG12ton259n83 );
splitter_AQFP splitterG13ton111n80_( clk_2 , G13 , 0 , splitterG13ton111n80 );
splitter_AQFP splitterG13ton262n80_( clk_3 , splitterG13ton111n80 , 0 , splitterG13ton262n80 );
splitter_AQFP splitterG14ton103n265_( clk_2 , G14 , 0 , splitterG14ton103n265 );
splitter_AQFP splitterG14ton181n265_( clk_5 , splitterG14ton103n265 , 0 , splitterG14ton181n265 );
splitter_AQFP splitterG15ton134n62_( clk_2 , G15 , 0 , splitterG15ton134n62 );
splitter_AQFP splitterG15ton227n62_( clk_3 , splitterG15ton134n62 , 0 , splitterG15ton227n62 );
splitter_AQFP splitterG16ton106n65_( clk_5 , buf_G16_splitterG16ton106n65_2 , 0 , splitterG16ton106n65 );
splitter_AQFP splitterG16ton230n65_( clk_6 , splitterG16ton106n65 , 0 , splitterG16ton230n65 );
splitter_AQFP splitterfromG17_( clk_4 , buf_G17_splitterfromG17_1 , 0 , splitterfromG17 );
splitter_AQFP splitterfromG18_( clk_5 , buf_G18_splitterfromG18_1 , 0 , splitterfromG18 );
splitter_AQFP splitterfromG19_( clk_6 , buf_G19_splitterfromG19_2 , 0 , splitterfromG19 );
splitter_AQFP splitterG2ton146n46_( clk_2 , G2 , 0 , splitterG2ton146n46 );
splitter_AQFP splitterG2ton211n46_( clk_3 , splitterG2ton146n46 , 0 , splitterG2ton211n46 );
splitter_AQFP splitterfromG20_( clk_4 , buf_G20_splitterfromG20_1 , 0 , splitterfromG20 );
splitter_AQFP splitterfromG21_( clk_3 , G21 , 0 , splitterfromG21 );
splitter_AQFP splitterfromG22_( clk_4 , buf_G22_splitterfromG22_1 , 0 , splitterfromG22 );
splitter_AQFP splitterG23ton109n200_( clk_3 , G23 , 0 , splitterG23ton109n200 );
splitter_AQFP splitterG24ton200n88_( clk_3 , buf_G24_splitterG24ton200n88_1 , 0 , splitterG24ton200n88 );
splitter_AQFP splitterG25ton193n281_( clk_3 , buf_G25_splitterG25ton193n281_9 , 0 , splitterG25ton193n281 );
splitter_AQFP splitterG26ton100n320_( clk_1 , buf_G26_splitterG26ton100n320_7 , 0 , splitterG26ton100n320 );
splitter_AQFP splitterG27ton153n287_( clk_1 , buf_G27_splitterG27ton153n287_7 , 0 , splitterG27ton153n287 );
splitter_AQFP splitterG28ton173n291_( clk_1 , buf_G28_splitterG28ton173n291_8 , 0 , splitterG28ton173n291 );
splitter_AQFP splitterfromG29_( clk_3 , buf_G29_splitterfromG29_1 , 0 , splitterfromG29 );
splitter_AQFP splitterG3ton156n46_( clk_2 , G3 , 0 , splitterG3ton156n46 );
splitter_AQFP splitterG3ton214n46_( clk_3 , splitterG3ton156n46 , 0 , splitterG3ton214n46 );
splitter_AQFP splitterfromG30_( clk_3 , buf_G30_splitterfromG30_1 , 0 , splitterfromG30 );
splitter_AQFP splitterG31ton126n99_( clk_2 , G31 , 0 , splitterG31ton126n99 );
splitter_AQFP splitterG31ton126n127_( clk_4 , splitterG31ton126n99 , 0 , splitterG31ton126n127 );
splitter_AQFP splitterG31ton152n201_( clk_5 , splitterG31ton126n99 , 0 , splitterG31ton152n201 );
splitter_AQFP splitterG31ton276n291_( clk_3 , splitterG31ton126n99 , 0 , splitterG31ton276n291 );
splitter_AQFP splitterG31ton295n99_( clk_2 , splitterG31ton126n99 , 0 , splitterG31ton295n99 );
splitter_AQFP splitterfromG32_( clk_6 , buf_G32_splitterfromG32_3 , 0 , splitterfromG32 );
splitter_AQFP splitterG33ton109n88_( clk_2 , G33 , 0 , splitterG33ton109n88 );
splitter_AQFP splitterG33ton199n273_( clk_4 , splitterG33ton109n88 , 0 , splitterG33ton199n273 );
splitter_AQFP splitterG33ton304n88_( clk_3 , splitterG33ton109n88 , 0 , splitterG33ton304n88 );
splitter_AQFP splitterG4ton117n43_( clk_2 , G4 , 0 , splitterG4ton117n43 );
splitter_AQFP splitterG4ton180n181_( clk_4 , splitterG4ton117n43 , 0 , splitterG4ton180n181 );
splitter_AQFP splitterG4ton216n43_( clk_6 , splitterG4ton117n43 , 0 , splitterG4ton216n43 );
splitter_AQFP splitterG5ton143n40_( clk_2 , G5 , 0 , splitterG5ton143n40 );
splitter_AQFP splitterG5ton237n40_( clk_7 , splitterG5ton143n40 , 0 , splitterG5ton237n40 );
splitter_AQFP splitterG6ton156n37_( clk_3 , G6 , 0 , splitterG6ton156n37 );
splitter_AQFP splitterG6ton240n37_( clk_4 , splitterG6ton156n37 , 0 , splitterG6ton240n37 );
splitter_AQFP splitterG7ton117n37_( clk_2 , G7 , 0 , splitterG7ton117n37 );
splitter_AQFP splitterG7ton243n37_( clk_4 , splitterG7ton117n37 , 0 , splitterG7ton243n37 );
splitter_AQFP splitterG8ton143n43_( clk_2 , G8 , 0 , splitterG8ton143n43 );
splitter_AQFP splitterG8ton159n160_( clk_1 , splitterG8ton143n43 , 0 , splitterG8ton159n160 );
splitter_AQFP splitterG8ton245n43_( clk_6 , splitterG8ton143n43 , 0 , splitterG8ton245n43 );
splitter_AQFP splitterG9ton103n59_( clk_3 , G9 , 0 , splitterG9ton103n59 );
splitter_AQFP splitterG9ton250n59_( clk_8 , splitterG9ton103n59 , 0 , splitterG9ton250n59 );
splitter_AQFP splitterfromn34_( clk_4 , n34 , 0 , splitterfromn34 );
splitter_AQFP splittern35ton252n78_( clk_4 , buf_n35_splittern35ton252n78_3 , 0 , splittern35ton252n78 );
splitter_AQFP splitterfromn38_( clk_7 , n38 , 0 , splitterfromn38 );
splitter_AQFP splittern41ton54n94_( clk_2 , n41 , 0 , splittern41ton54n94 );
splitter_AQFP splitterfromn44_( clk_1 , n44 , 0 , splitterfromn44 );
splitter_AQFP splitterfromn47_( clk_6 , n47 , 0 , splitterfromn47 );
splitter_AQFP splittern50ton186n52_( clk_1 , n50 , 0 , splittern50ton186n52 );
splitter_AQFP splitterfromn53_( clk_4 , n53 , 0 , splitterfromn53 );
splitter_AQFP splittern56ton299n71_( clk_7 , n56 , 0 , splittern56ton299n71 );
splitter_AQFP splitterfromn57_( clk_8 , buf_n57_splitterfromn57_1 , 0 , splitterfromn57 );
splitter_AQFP splitterfromn60_( clk_3 , n60 , 0 , splitterfromn60 );
splitter_AQFP splittern63ton163n65_( clk_6 , n63 , 0 , splittern63ton163n65 );
splitter_AQFP splittern66ton67n86_( clk_1 , n66 , 0 , splittern66ton67n86 );
splitter_AQFP splitterfromn69_( clk_7 , n69 , 0 , splitterfromn69 );
splitter_AQFP splitterfromn72_( clk_2 , n72 , 0 , splitterfromn72 );
splitter_AQFP splittern73ton278n76_( clk_4 , n73 , 0 , splittern73ton278n76 );
splitter_AQFP splittern74ton275n76_( clk_3 , buf_n74_splittern74ton275n76_1 , 0 , splittern74ton275n76 );
splitter_AQFP splittern77ton253n78_( clk_7 , n77 , 0 , splittern77ton253n78 );
splitter_AQFP splitterfromn78_( clk_1 , n78 , 0 , splitterfromn78 );
splitter_AQFP splitterfromn81_( clk_6 , n81 , 0 , splitterfromn81 );
splitter_AQFP splitterfromn84_( clk_1 , n84 , 0 , splitterfromn84 );
splitter_AQFP splittern87ton189n97_( clk_4 , n87 , 0 , splittern87ton189n97 );
splitter_AQFP splittern87ton309n97_( clk_5 , splittern87ton189n97 , 0 , splittern87ton309n97 );
splitter_AQFP splitterfromn88_( clk_5 , n88 , 0 , splitterfromn88 );
splitter_AQFP splitterfromn89_( clk_7 , n89 , 0 , splitterfromn89 );
splitter_AQFP splitterfromn92_( clk_2 , n92 , 0 , splitterfromn92 );
splitter_AQFP splitterfromn95_( clk_5 , n95 , 0 , splitterfromn95 );
splitter_AQFP splitterfromn98_( clk_8 , n98 , 0 , splitterfromn98 );
splitter_AQFP splitterfromn99_( clk_2 , n99 , 0 , splitterfromn99 );
splitter_AQFP splittern105ton106n309_( clk_6 , n105 , 0 , splittern105ton106n309 );
splitter_AQFP splittern108ton114n141_( clk_2 , n108 , 0 , splittern108ton114n141 );
splitter_AQFP splitterfromn109_( clk_5 , n109 , 0 , splitterfromn109 );
splitter_AQFP splitterfromn110_( clk_7 , n110 , 0 , splitterfromn110 );
splitter_AQFP splitterfromn113_( clk_2 , n113 , 0 , splitterfromn113 );
splitter_AQFP splitterfromn116_( clk_5 , n116 , 0 , splitterfromn116 );
splitter_AQFP splitterfromn119_( clk_5 , n119 , 0 , splitterfromn119 );
splitter_AQFP splitterfromn122_( clk_4 , buf_n122_splitterfromn122_1 , 0 , splitterfromn122 );
splitter_AQFP splitterfromn125_( clk_8 , n125 , 0 , splitterfromn125 );
splitter_AQFP splitterfromn126_( clk_2 , n126 , 0 , splitterfromn126 );
splitter_AQFP splitterfromn127_( clk_7 , n127 , 0 , splitterfromn127 );
splitter_AQFP splittern128ton129n295_( clk_2 , n128 , 0 , splittern128ton129n295 );
splitter_AQFP splitterfromn133_( clk_7 , n133 , 0 , splitterfromn133 );
splitter_AQFP splitterfromn136_( clk_6 , n136 , 0 , splitterfromn136 );
splitter_AQFP splitterfromn139_( clk_2 , n139 , 0 , splitterfromn139 );
splitter_AQFP splitterfromn142_( clk_5 , n142 , 0 , splitterfromn142 );
splitter_AQFP splitterfromn145_( clk_5 , n145 , 0 , splitterfromn145 );
splitter_AQFP splitterfromn148_( clk_4 , buf_n148_splitterfromn148_2 , 0 , splitterfromn148 );
splitter_AQFP splitterfromn151_( clk_8 , n151 , 0 , splitterfromn151 );
splitter_AQFP splitterfromn152_( clk_2 , n152 , 0 , splitterfromn152 );
splitter_AQFP splitterfromn158_( clk_8 , n158 , 0 , splitterfromn158 );
splitter_AQFP splitterfromn161_( clk_4 , n161 , 0 , splitterfromn161 );
splitter_AQFP splitterfromn162_( clk_8 , n162 , 0 , splitterfromn162 );
splitter_AQFP splitterfromn165_( clk_1 , n165 , 0 , splitterfromn165 );
splitter_AQFP splitterfromn168_( clk_4 , n168 , 0 , splitterfromn168 );
splitter_AQFP splitterfromn171_( clk_8 , n171 , 0 , splitterfromn171 );
splitter_AQFP splitterfromn172_( clk_2 , n172 , 0 , splitterfromn172 );
splitter_AQFP splittern177ton197n272_( clk_7 , n177 , 0 , splittern177ton197n272 );
splitter_AQFP splittern178ton196n269_( clk_5 , buf_n178_splittern178ton196n269_2 , 0 , splittern178ton196n269 );
splitter_AQFP splitterfromn179_( clk_7 , n179 , 0 , splitterfromn179 );
splitter_AQFP splitterfromn182_( clk_8 , n182 , 0 , splitterfromn182 );
splitter_AQFP splitterfromn185_( clk_3 , n185 , 0 , splitterfromn185 );
splitter_AQFP splitterfromn188_( clk_6 , n188 , 0 , splitterfromn188 );
splitter_AQFP splitterfromn191_( clk_1 , n191 , 0 , splitterfromn191 );
splitter_AQFP splittern192ton193n284_( clk_3 , n192 , 0 , splittern192ton193n284 );
splitter_AQFP splittern195ton196n270_( clk_6 , n195 , 0 , splittern195ton196n270 );
splitter_AQFP splitterfromn197_( clk_1 , n197 , 0 , splitterfromn197 );
splitter_AQFP splitterfromn198_( clk_3 , n198 , 0 , splitterfromn198 );
splitter_AQFP splitterfromn199_( clk_6 , buf_n199_splitterfromn199_3 , 0 , splitterfromn199 );
splitter_AQFP splitterfromn200_( clk_4 , buf_n200_splitterfromn200_2 , 0 , splitterfromn200 );
splitter_AQFP splitterfromn201_( clk_7 , n201 , 0 , splitterfromn201 );
splitter_AQFP splittern203ton204n321_( clk_6 , buf_n203_splittern203ton204n321_3 , 0 , splittern203ton204n321 );
splitter_AQFP splittern203ton290n321_( clk_2 , splittern203ton204n321 , 0 , splittern203ton290n321 );
splitter_AQFP splitterfromn204_( clk_1 , n204 , 0 , splitterfromn204 );
splitter_AQFP splitterfromn205_( clk_4 , n205 , 0 , splitterfromn205 );
splitter_AQFP splittern206ton207n302_( clk_5 , n206 , 0 , splittern206ton207n302 );
splitter_AQFP splittern206ton208n210_( clk_6 , splittern206ton207n302 , 0 , splittern206ton208n210 );
splitter_AQFP splittern206ton211n216_( clk_6 , splittern206ton207n302 , 0 , splittern206ton211n216 );
splitter_AQFP splittern206ton217n302_( clk_6 , splittern206ton207n302 , 0 , splittern206ton217n302 );
splitter_AQFP splitterfromn219_( clk_7 , buf_n219_splitterfromn219_5 , 0 , splitterfromn219 );
splitter_AQFP splittern221ton222n254_( clk_7 , buf_n221_splittern221ton222n254_2 , 0 , splittern221ton222n254 );
splitter_AQFP splittern222ton223n314_( clk_5 , n222 , 0 , splittern222ton223n314 );
splitter_AQFP splittern222ton226n229_( clk_6 , splittern222ton223n314 , 0 , splittern222ton226n229 );
splitter_AQFP splittern222ton230n314_( clk_6 , splittern222ton223n314 , 0 , splittern222ton230n314 );
splitter_AQFP splitterfromn234_( clk_3 , n234 , 0 , splitterfromn234 );
splitter_AQFP splittern235ton236n246_( clk_5 , n235 , 0 , splittern235ton236n246 );
splitter_AQFP splittern235ton239n240_( clk_6 , splittern235ton236n246 , 0 , splittern235ton239n240 );
splitter_AQFP splittern235ton242n246_( clk_6 , splittern235ton236n246 , 0 , splittern235ton242n246 );
splitter_AQFP splitterfromn248_( clk_5 , n248 , 0 , splitterfromn248 );
splitter_AQFP splittern254ton255n265_( clk_5 , n254 , 0 , splittern254ton255n265 );
splitter_AQFP splittern254ton258n259_( clk_6 , splittern254ton255n265 , 0 , splittern254ton258n259 );
splitter_AQFP splittern254ton261n265_( clk_6 , splittern254ton255n265 , 0 , splittern254ton261n265 );
splitter_AQFP splittern267ton268n320_( clk_8 , n267 , 0 , splittern267ton268n320 );
splitter_AQFP splittern267ton288n320_( clk_1 , splittern267ton268n320 , 0 , splittern267ton288n320 );
splitter_AQFP splitterfromn275_( clk_2 , n275 , 0 , splitterfromn275 );
splitter_AQFP splitterfromn281_( clk_2 , n281 , 0 , splitterfromn281 );
splitter_AQFP splitterfromn299_( clk_1 , n299 , 0 , splitterfromn299 );
splitter_AQFP splitterfromn300_( clk_6 , buf_n300_splitterfromn300_5 , 0 , splitterfromn300 );
splitter_AQFP splitterfromn304_( clk_2 , n304 , 0 , splitterfromn304 );
splitter_AQFP splitterfromn311_( clk_3 , buf_n311_splitterfromn311_3 , 0 , splitterfromn311 );
splitter_AQFP splitterfromn312_( clk_5 , buf_n312_splitterfromn312_4 , 0 , splitterfromn312 );
splitter_AQFP splitterfromn316_( clk_2 , n316 , 0 , splitterfromn316 );

endmodule