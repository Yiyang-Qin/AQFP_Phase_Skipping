module top( clk_1 , clk_2 , clk_3 , clk_4 , clk_5 , clk_6 , clk_7 , clk_8 , G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G5 , G6 , G7 , G8 , G9 , G1324 , G1325 , G1326 , G1327 , G1328 , G1329 , G1330 , G1331 , G1332 , G1333 , G1334 , G1335 , G1336 , G1337 , G1338 , G1339 , G1340 , G1341 , G1342 , G1343 , G1344 , G1345 , G1346 , G1347 , G1348 , G1349 , G1350 , G1351 , G1352 , G1353 , G1354 , G1355 );

input G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G5 , G6 , G7 , G8 , G9 ;
output G1324 , G1325 , G1326 , G1327 , G1328 , G1329 , G1330 , G1331 , G1332 , G1333 , G1334 , G1335 , G1336 , G1337 , G1338 , G1339 , G1340 , G1341 , G1342 , G1343 , G1344 , G1345 , G1346 , G1347 , G1348 , G1349 , G1350 , G1351 , G1352 , G1353 , G1354 , G1355 ;
wire n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , buf_G33_n42_1 , buf_G34_n193_1 , buf_G35_n231_1 , buf_G36_n254_1 , buf_G37_n154_1 , buf_G39_n88_1 , buf_G40_n125_1 , buf_n42_splitterfromn42_1 , buf_n88_splitterfromn88_1 , buf_n125_splitterfromn125_1 , buf_n154_splitterfromn154_1 , buf_n173_splitterfromn173_2 , buf_n173_splitterfromn173_1 , buf_n193_splitterfromn193_1 , buf_n231_splitterfromn231_1 , buf_n254_splitterfromn254_1 , buf_n383_G1344_1 , buf_n387_G1345_1 , buf_n391_G1346_1 , buf_n395_G1347_1 , buf_n418_G1352_1 , buf_n422_G1353_1 , buf_n426_G1354_1 , buf_n430_G1355_1 , buf_splitterG1ton83n284_splitterG1ton283n284_12 , buf_splitterG1ton83n284_splitterG1ton283n284_11 , buf_splitterG1ton83n284_splitterG1ton283n284_10 , buf_splitterG1ton83n284_splitterG1ton283n284_9 , buf_splitterG1ton83n284_splitterG1ton283n284_8 , buf_splitterG1ton83n284_splitterG1ton283n284_7 , buf_splitterG1ton83n284_splitterG1ton283n284_6 , buf_splitterG1ton83n284_splitterG1ton283n284_5 , buf_splitterG1ton83n284_splitterG1ton283n284_4 , buf_splitterG1ton83n284_splitterG1ton283n284_3 , buf_splitterG1ton83n284_splitterG1ton283n284_2 , buf_splitterG1ton83n284_splitterG1ton283n284_1 , buf_splitterG10ton219n325_splitterG10ton324n325_11 , buf_splitterG10ton219n325_splitterG10ton324n325_10 , buf_splitterG10ton219n325_splitterG10ton324n325_9 , buf_splitterG10ton219n325_splitterG10ton324n325_8 , buf_splitterG10ton219n325_splitterG10ton324n325_7 , buf_splitterG10ton219n325_splitterG10ton324n325_6 , buf_splitterG10ton219n325_splitterG10ton324n325_5 , buf_splitterG10ton219n325_splitterG10ton324n325_4 , buf_splitterG10ton219n325_splitterG10ton324n325_3 , buf_splitterG10ton219n325_splitterG10ton324n325_2 , buf_splitterG10ton219n325_splitterG10ton324n325_1 , buf_splitterG11ton235n329_splitterG11ton328n329_11 , buf_splitterG11ton235n329_splitterG11ton328n329_10 , buf_splitterG11ton235n329_splitterG11ton328n329_9 , buf_splitterG11ton235n329_splitterG11ton328n329_8 , buf_splitterG11ton235n329_splitterG11ton328n329_7 , buf_splitterG11ton235n329_splitterG11ton328n329_6 , buf_splitterG11ton235n329_splitterG11ton328n329_5 , buf_splitterG11ton235n329_splitterG11ton328n329_4 , buf_splitterG11ton235n329_splitterG11ton328n329_3 , buf_splitterG11ton235n329_splitterG11ton328n329_2 , buf_splitterG11ton235n329_splitterG11ton328n329_1 , buf_splitterG12ton93n333_splitterG12ton332n333_11 , buf_splitterG12ton93n333_splitterG12ton332n333_10 , buf_splitterG12ton93n333_splitterG12ton332n333_9 , buf_splitterG12ton93n333_splitterG12ton332n333_8 , buf_splitterG12ton93n333_splitterG12ton332n333_7 , buf_splitterG12ton93n333_splitterG12ton332n333_6 , buf_splitterG12ton93n333_splitterG12ton332n333_5 , buf_splitterG12ton93n333_splitterG12ton332n333_4 , buf_splitterG12ton93n333_splitterG12ton332n333_3 , buf_splitterG12ton93n333_splitterG12ton332n333_2 , buf_splitterG12ton93n333_splitterG12ton332n333_1 , buf_splitterG13ton65n339_splitterG13ton338n339_11 , buf_splitterG13ton65n339_splitterG13ton338n339_10 , buf_splitterG13ton65n339_splitterG13ton338n339_9 , buf_splitterG13ton65n339_splitterG13ton338n339_8 , buf_splitterG13ton65n339_splitterG13ton338n339_7 , buf_splitterG13ton65n339_splitterG13ton338n339_6 , buf_splitterG13ton65n339_splitterG13ton338n339_5 , buf_splitterG13ton65n339_splitterG13ton338n339_4 , buf_splitterG13ton65n339_splitterG13ton338n339_3 , buf_splitterG13ton65n339_splitterG13ton338n339_2 , buf_splitterG13ton65n339_splitterG13ton338n339_1 , buf_splitterG14ton216n343_splitterG14ton342n343_11 , buf_splitterG14ton216n343_splitterG14ton342n343_10 , buf_splitterG14ton216n343_splitterG14ton342n343_9 , buf_splitterG14ton216n343_splitterG14ton342n343_8 , buf_splitterG14ton216n343_splitterG14ton342n343_7 , buf_splitterG14ton216n343_splitterG14ton342n343_6 , buf_splitterG14ton216n343_splitterG14ton342n343_5 , buf_splitterG14ton216n343_splitterG14ton342n343_4 , buf_splitterG14ton216n343_splitterG14ton342n343_3 , buf_splitterG14ton216n343_splitterG14ton342n343_2 , buf_splitterG14ton216n343_splitterG14ton342n343_1 , buf_splitterG15ton236n347_splitterG15ton346n347_10 , buf_splitterG15ton236n347_splitterG15ton346n347_9 , buf_splitterG15ton236n347_splitterG15ton346n347_8 , buf_splitterG15ton236n347_splitterG15ton346n347_7 , buf_splitterG15ton236n347_splitterG15ton346n347_6 , buf_splitterG15ton236n347_splitterG15ton346n347_5 , buf_splitterG15ton236n347_splitterG15ton346n347_4 , buf_splitterG15ton236n347_splitterG15ton346n347_3 , buf_splitterG15ton236n347_splitterG15ton346n347_2 , buf_splitterG15ton236n347_splitterG15ton346n347_1 , buf_splitterG16ton262n351_splitterG16ton350n351_10 , buf_splitterG16ton262n351_splitterG16ton350n351_9 , buf_splitterG16ton262n351_splitterG16ton350n351_8 , buf_splitterG16ton262n351_splitterG16ton350n351_7 , buf_splitterG16ton262n351_splitterG16ton350n351_6 , buf_splitterG16ton262n351_splitterG16ton350n351_5 , buf_splitterG16ton262n351_splitterG16ton350n351_4 , buf_splitterG16ton262n351_splitterG16ton350n351_3 , buf_splitterG16ton262n351_splitterG16ton350n351_2 , buf_splitterG16ton262n351_splitterG16ton350n351_1 , buf_splitterG17ton44n364_splitterG17ton363n364_11 , buf_splitterG17ton44n364_splitterG17ton363n364_10 , buf_splitterG17ton44n364_splitterG17ton363n364_9 , buf_splitterG17ton44n364_splitterG17ton363n364_8 , buf_splitterG17ton44n364_splitterG17ton363n364_7 , buf_splitterG17ton44n364_splitterG17ton363n364_6 , buf_splitterG17ton44n364_splitterG17ton363n364_5 , buf_splitterG17ton44n364_splitterG17ton363n364_4 , buf_splitterG17ton44n364_splitterG17ton363n364_3 , buf_splitterG17ton44n364_splitterG17ton363n364_2 , buf_splitterG17ton44n364_splitterG17ton363n364_1 , buf_splitterG18ton47n368_splitterG18ton367n368_11 , buf_splitterG18ton47n368_splitterG18ton367n368_10 , buf_splitterG18ton47n368_splitterG18ton367n368_9 , buf_splitterG18ton47n368_splitterG18ton367n368_8 , buf_splitterG18ton47n368_splitterG18ton367n368_7 , buf_splitterG18ton47n368_splitterG18ton367n368_6 , buf_splitterG18ton47n368_splitterG18ton367n368_5 , buf_splitterG18ton47n368_splitterG18ton367n368_4 , buf_splitterG18ton47n368_splitterG18ton367n368_3 , buf_splitterG18ton47n368_splitterG18ton367n368_2 , buf_splitterG18ton47n368_splitterG18ton367n368_1 , buf_splitterG19ton44n372_splitterG19ton371n372_11 , buf_splitterG19ton44n372_splitterG19ton371n372_10 , buf_splitterG19ton44n372_splitterG19ton371n372_9 , buf_splitterG19ton44n372_splitterG19ton371n372_8 , buf_splitterG19ton44n372_splitterG19ton371n372_7 , buf_splitterG19ton44n372_splitterG19ton371n372_6 , buf_splitterG19ton44n372_splitterG19ton371n372_5 , buf_splitterG19ton44n372_splitterG19ton371n372_4 , buf_splitterG19ton44n372_splitterG19ton371n372_3 , buf_splitterG19ton44n372_splitterG19ton371n372_2 , buf_splitterG19ton44n372_splitterG19ton371n372_1 , buf_splitterG2ton216n288_splitterG2ton287n288_12 , buf_splitterG2ton216n288_splitterG2ton287n288_11 , buf_splitterG2ton216n288_splitterG2ton287n288_10 , buf_splitterG2ton216n288_splitterG2ton287n288_9 , buf_splitterG2ton216n288_splitterG2ton287n288_8 , buf_splitterG2ton216n288_splitterG2ton287n288_7 , buf_splitterG2ton216n288_splitterG2ton287n288_6 , buf_splitterG2ton216n288_splitterG2ton287n288_5 , buf_splitterG2ton216n288_splitterG2ton287n288_4 , buf_splitterG2ton216n288_splitterG2ton287n288_3 , buf_splitterG2ton216n288_splitterG2ton287n288_2 , buf_splitterG2ton216n288_splitterG2ton287n288_1 , buf_splitterG20ton47n376_splitterG20ton375n376_11 , buf_splitterG20ton47n376_splitterG20ton375n376_10 , buf_splitterG20ton47n376_splitterG20ton375n376_9 , buf_splitterG20ton47n376_splitterG20ton375n376_8 , buf_splitterG20ton47n376_splitterG20ton375n376_7 , buf_splitterG20ton47n376_splitterG20ton375n376_6 , buf_splitterG20ton47n376_splitterG20ton375n376_5 , buf_splitterG20ton47n376_splitterG20ton375n376_4 , buf_splitterG20ton47n376_splitterG20ton375n376_3 , buf_splitterG20ton47n376_splitterG20ton375n376_2 , buf_splitterG20ton47n376_splitterG20ton375n376_1 , buf_splitterG21ton59n382_splitterG21ton381n382_10 , buf_splitterG21ton59n382_splitterG21ton381n382_9 , buf_splitterG21ton59n382_splitterG21ton381n382_8 , buf_splitterG21ton59n382_splitterG21ton381n382_7 , buf_splitterG21ton59n382_splitterG21ton381n382_6 , buf_splitterG21ton59n382_splitterG21ton381n382_5 , buf_splitterG21ton59n382_splitterG21ton381n382_4 , buf_splitterG21ton59n382_splitterG21ton381n382_3 , buf_splitterG21ton59n382_splitterG21ton381n382_2 , buf_splitterG21ton59n382_splitterG21ton381n382_1 , buf_splitterG22ton56n386_splitterG22ton385n386_10 , buf_splitterG22ton56n386_splitterG22ton385n386_9 , buf_splitterG22ton56n386_splitterG22ton385n386_8 , buf_splitterG22ton56n386_splitterG22ton385n386_7 , buf_splitterG22ton56n386_splitterG22ton385n386_6 , buf_splitterG22ton56n386_splitterG22ton385n386_5 , buf_splitterG22ton56n386_splitterG22ton385n386_4 , buf_splitterG22ton56n386_splitterG22ton385n386_3 , buf_splitterG22ton56n386_splitterG22ton385n386_2 , buf_splitterG22ton56n386_splitterG22ton385n386_1 , buf_splitterG23ton56n390_splitterG23ton389n390_10 , buf_splitterG23ton56n390_splitterG23ton389n390_9 , buf_splitterG23ton56n390_splitterG23ton389n390_8 , buf_splitterG23ton56n390_splitterG23ton389n390_7 , buf_splitterG23ton56n390_splitterG23ton389n390_6 , buf_splitterG23ton56n390_splitterG23ton389n390_5 , buf_splitterG23ton56n390_splitterG23ton389n390_4 , buf_splitterG23ton56n390_splitterG23ton389n390_3 , buf_splitterG23ton56n390_splitterG23ton389n390_2 , buf_splitterG23ton56n390_splitterG23ton389n390_1 , buf_splitterG24ton59n394_splitterG24ton393n394_10 , buf_splitterG24ton59n394_splitterG24ton393n394_9 , buf_splitterG24ton59n394_splitterG24ton393n394_8 , buf_splitterG24ton59n394_splitterG24ton393n394_7 , buf_splitterG24ton59n394_splitterG24ton393n394_6 , buf_splitterG24ton59n394_splitterG24ton393n394_5 , buf_splitterG24ton59n394_splitterG24ton393n394_4 , buf_splitterG24ton59n394_splitterG24ton393n394_3 , buf_splitterG24ton59n394_splitterG24ton393n394_2 , buf_splitterG24ton59n394_splitterG24ton393n394_1 , buf_splitterG25ton207n399_splitterG25ton398n399_11 , buf_splitterG25ton207n399_splitterG25ton398n399_10 , buf_splitterG25ton207n399_splitterG25ton398n399_9 , buf_splitterG25ton207n399_splitterG25ton398n399_8 , buf_splitterG25ton207n399_splitterG25ton398n399_7 , buf_splitterG25ton207n399_splitterG25ton398n399_6 , buf_splitterG25ton207n399_splitterG25ton398n399_5 , buf_splitterG25ton207n399_splitterG25ton398n399_4 , buf_splitterG25ton207n399_splitterG25ton398n399_3 , buf_splitterG25ton207n399_splitterG25ton398n399_2 , buf_splitterG25ton207n399_splitterG25ton398n399_1 , buf_splitterG26ton210n403_splitterG26ton402n403_11 , buf_splitterG26ton210n403_splitterG26ton402n403_10 , buf_splitterG26ton210n403_splitterG26ton402n403_9 , buf_splitterG26ton210n403_splitterG26ton402n403_8 , buf_splitterG26ton210n403_splitterG26ton402n403_7 , buf_splitterG26ton210n403_splitterG26ton402n403_6 , buf_splitterG26ton210n403_splitterG26ton402n403_5 , buf_splitterG26ton210n403_splitterG26ton402n403_4 , buf_splitterG26ton210n403_splitterG26ton402n403_3 , buf_splitterG26ton210n403_splitterG26ton402n403_2 , buf_splitterG26ton210n403_splitterG26ton402n403_1 , buf_splitterG27ton210n407_splitterG27ton406n407_11 , buf_splitterG27ton210n407_splitterG27ton406n407_10 , buf_splitterG27ton210n407_splitterG27ton406n407_9 , buf_splitterG27ton210n407_splitterG27ton406n407_8 , buf_splitterG27ton210n407_splitterG27ton406n407_7 , buf_splitterG27ton210n407_splitterG27ton406n407_6 , buf_splitterG27ton210n407_splitterG27ton406n407_5 , buf_splitterG27ton210n407_splitterG27ton406n407_4 , buf_splitterG27ton210n407_splitterG27ton406n407_3 , buf_splitterG27ton210n407_splitterG27ton406n407_2 , buf_splitterG27ton210n407_splitterG27ton406n407_1 , buf_splitterG28ton207n411_splitterG28ton410n411_11 , buf_splitterG28ton207n411_splitterG28ton410n411_10 , buf_splitterG28ton207n411_splitterG28ton410n411_9 , buf_splitterG28ton207n411_splitterG28ton410n411_8 , buf_splitterG28ton207n411_splitterG28ton410n411_7 , buf_splitterG28ton207n411_splitterG28ton410n411_6 , buf_splitterG28ton207n411_splitterG28ton410n411_5 , buf_splitterG28ton207n411_splitterG28ton410n411_4 , buf_splitterG28ton207n411_splitterG28ton410n411_3 , buf_splitterG28ton207n411_splitterG28ton410n411_2 , buf_splitterG28ton207n411_splitterG28ton410n411_1 , buf_splitterG29ton195n417_splitterG29ton416n417_10 , buf_splitterG29ton195n417_splitterG29ton416n417_9 , buf_splitterG29ton195n417_splitterG29ton416n417_8 , buf_splitterG29ton195n417_splitterG29ton416n417_7 , buf_splitterG29ton195n417_splitterG29ton416n417_6 , buf_splitterG29ton195n417_splitterG29ton416n417_5 , buf_splitterG29ton195n417_splitterG29ton416n417_4 , buf_splitterG29ton195n417_splitterG29ton416n417_3 , buf_splitterG29ton195n417_splitterG29ton416n417_2 , buf_splitterG29ton195n417_splitterG29ton416n417_1 , buf_splitterG3ton239n292_splitterG3ton291n292_11 , buf_splitterG3ton239n292_splitterG3ton291n292_10 , buf_splitterG3ton239n292_splitterG3ton291n292_9 , buf_splitterG3ton239n292_splitterG3ton291n292_8 , buf_splitterG3ton239n292_splitterG3ton291n292_7 , buf_splitterG3ton239n292_splitterG3ton291n292_6 , buf_splitterG3ton239n292_splitterG3ton291n292_5 , buf_splitterG3ton239n292_splitterG3ton291n292_4 , buf_splitterG3ton239n292_splitterG3ton291n292_3 , buf_splitterG3ton239n292_splitterG3ton291n292_2 , buf_splitterG3ton239n292_splitterG3ton291n292_1 , buf_splitterG30ton195n421_splitterG30ton420n421_10 , buf_splitterG30ton195n421_splitterG30ton420n421_9 , buf_splitterG30ton195n421_splitterG30ton420n421_8 , buf_splitterG30ton195n421_splitterG30ton420n421_7 , buf_splitterG30ton195n421_splitterG30ton420n421_6 , buf_splitterG30ton195n421_splitterG30ton420n421_5 , buf_splitterG30ton195n421_splitterG30ton420n421_4 , buf_splitterG30ton195n421_splitterG30ton420n421_3 , buf_splitterG30ton195n421_splitterG30ton420n421_2 , buf_splitterG30ton195n421_splitterG30ton420n421_1 , buf_splitterG31ton198n425_splitterG31ton424n425_10 , buf_splitterG31ton198n425_splitterG31ton424n425_9 , buf_splitterG31ton198n425_splitterG31ton424n425_8 , buf_splitterG31ton198n425_splitterG31ton424n425_7 , buf_splitterG31ton198n425_splitterG31ton424n425_6 , buf_splitterG31ton198n425_splitterG31ton424n425_5 , buf_splitterG31ton198n425_splitterG31ton424n425_4 , buf_splitterG31ton198n425_splitterG31ton424n425_3 , buf_splitterG31ton198n425_splitterG31ton424n425_2 , buf_splitterG31ton198n425_splitterG31ton424n425_1 , buf_splitterG32ton198n429_splitterG32ton428n429_10 , buf_splitterG32ton198n429_splitterG32ton428n429_9 , buf_splitterG32ton198n429_splitterG32ton428n429_8 , buf_splitterG32ton198n429_splitterG32ton428n429_7 , buf_splitterG32ton198n429_splitterG32ton428n429_6 , buf_splitterG32ton198n429_splitterG32ton428n429_5 , buf_splitterG32ton198n429_splitterG32ton428n429_4 , buf_splitterG32ton198n429_splitterG32ton428n429_3 , buf_splitterG32ton198n429_splitterG32ton428n429_2 , buf_splitterG32ton198n429_splitterG32ton428n429_1 , buf_splitterG4ton80n296_splitterG4ton295n296_12 , buf_splitterG4ton80n296_splitterG4ton295n296_11 , buf_splitterG4ton80n296_splitterG4ton295n296_10 , buf_splitterG4ton80n296_splitterG4ton295n296_9 , buf_splitterG4ton80n296_splitterG4ton295n296_8 , buf_splitterG4ton80n296_splitterG4ton295n296_7 , buf_splitterG4ton80n296_splitterG4ton295n296_6 , buf_splitterG4ton80n296_splitterG4ton295n296_5 , buf_splitterG4ton80n296_splitterG4ton295n296_4 , buf_splitterG4ton80n296_splitterG4ton295n296_3 , buf_splitterG4ton80n296_splitterG4ton295n296_2 , buf_splitterG4ton80n296_splitterG4ton295n296_1 , buf_splitterG5ton65n302_splitterG5ton301n302_12 , buf_splitterG5ton65n302_splitterG5ton301n302_11 , buf_splitterG5ton65n302_splitterG5ton301n302_10 , buf_splitterG5ton65n302_splitterG5ton301n302_9 , buf_splitterG5ton65n302_splitterG5ton301n302_8 , buf_splitterG5ton65n302_splitterG5ton301n302_7 , buf_splitterG5ton65n302_splitterG5ton301n302_6 , buf_splitterG5ton65n302_splitterG5ton301n302_5 , buf_splitterG5ton65n302_splitterG5ton301n302_4 , buf_splitterG5ton65n302_splitterG5ton301n302_3 , buf_splitterG5ton65n302_splitterG5ton301n302_2 , buf_splitterG5ton65n302_splitterG5ton301n302_1 , buf_splitterG6ton219n306_splitterG6ton305n306_12 , buf_splitterG6ton219n306_splitterG6ton305n306_11 , buf_splitterG6ton219n306_splitterG6ton305n306_10 , buf_splitterG6ton219n306_splitterG6ton305n306_9 , buf_splitterG6ton219n306_splitterG6ton305n306_8 , buf_splitterG6ton219n306_splitterG6ton305n306_7 , buf_splitterG6ton219n306_splitterG6ton305n306_6 , buf_splitterG6ton219n306_splitterG6ton305n306_5 , buf_splitterG6ton219n306_splitterG6ton305n306_4 , buf_splitterG6ton219n306_splitterG6ton305n306_3 , buf_splitterG6ton219n306_splitterG6ton305n306_2 , buf_splitterG6ton219n306_splitterG6ton305n306_1 , buf_splitterG7ton239n310_splitterG7ton309n310_11 , buf_splitterG7ton239n310_splitterG7ton309n310_10 , buf_splitterG7ton239n310_splitterG7ton309n310_9 , buf_splitterG7ton239n310_splitterG7ton309n310_8 , buf_splitterG7ton239n310_splitterG7ton309n310_7 , buf_splitterG7ton239n310_splitterG7ton309n310_6 , buf_splitterG7ton239n310_splitterG7ton309n310_5 , buf_splitterG7ton239n310_splitterG7ton309n310_4 , buf_splitterG7ton239n310_splitterG7ton309n310_3 , buf_splitterG7ton239n310_splitterG7ton309n310_2 , buf_splitterG7ton239n310_splitterG7ton309n310_1 , buf_splitterG8ton262n314_splitterG8ton313n314_11 , buf_splitterG8ton262n314_splitterG8ton313n314_10 , buf_splitterG8ton262n314_splitterG8ton313n314_9 , buf_splitterG8ton262n314_splitterG8ton313n314_8 , buf_splitterG8ton262n314_splitterG8ton313n314_7 , buf_splitterG8ton262n314_splitterG8ton313n314_6 , buf_splitterG8ton262n314_splitterG8ton313n314_5 , buf_splitterG8ton262n314_splitterG8ton313n314_4 , buf_splitterG8ton262n314_splitterG8ton313n314_3 , buf_splitterG8ton262n314_splitterG8ton313n314_2 , buf_splitterG8ton262n314_splitterG8ton313n314_1 , buf_splitterG9ton96n321_splitterG9ton320n321_11 , buf_splitterG9ton96n321_splitterG9ton320n321_10 , buf_splitterG9ton96n321_splitterG9ton320n321_9 , buf_splitterG9ton96n321_splitterG9ton320n321_8 , buf_splitterG9ton96n321_splitterG9ton320n321_7 , buf_splitterG9ton96n321_splitterG9ton320n321_6 , buf_splitterG9ton96n321_splitterG9ton320n321_5 , buf_splitterG9ton96n321_splitterG9ton320n321_4 , buf_splitterG9ton96n321_splitterG9ton320n321_3 , buf_splitterG9ton96n321_splitterG9ton320n321_2 , buf_splitterG9ton96n321_splitterG9ton320n321_1 , buf_splittern78ton230n300_splittern78ton277n300_1 , buf_splittern78ton277n300_splittern78ton337n300_2 , buf_splittern78ton277n300_splittern78ton337n300_1 , buf_splittern115ton354n405_splittern115ton388n405_2 , buf_splittern115ton354n405_splittern115ton388n405_1 , buf_splittern152ton354n409_splittern152ton392n409_2 , buf_splittern152ton354n409_splittern152ton392n409_1 , buf_splittern153ton356n281_splittern153ton317n281_2 , buf_splittern153ton356n281_splittern153ton317n281_1 , buf_splittern153ton317n281_n281_1 , buf_splittern172ton357n397_splittern172ton380n397_2 , buf_splittern172ton357n397_splittern172ton380n397_1 , buf_splittern191ton357n401_splittern191ton384n401_2 , buf_splittern191ton357n401_splittern191ton384n401_1 , buf_splitterfromn192_n280_3 , buf_splitterfromn192_n280_2 , buf_splitterfromn192_n280_1 , buf_splittern229ton277n304_splittern229ton341n304_3 , buf_splittern229ton277n304_splittern229ton341n304_2 , buf_splittern229ton277n304_splittern229ton341n304_1 , buf_splitterfromn230_n396_3 , buf_splitterfromn230_n396_2 , buf_splitterfromn230_n396_1 , buf_splittern249ton275n308_splittern249ton345n308_2 , buf_splittern249ton275n308_splittern249ton345n308_1 , buf_splitterfromn251_n361_3 , buf_splitterfromn251_n361_2 , buf_splitterfromn251_n361_1 , buf_splittern272ton273n312_splittern272ton349n312_1 , buf_splitterfromn274_n360_1 , buf_splittern298ton356n299_splittern298ton335n299_1 , buf_splittern298ton335n299_n299_2 , buf_splittern298ton335n299_n299_1 , buf_splittern316ton353n318_splittern316ton335n318_1 , buf_splittern316ton335n318_n318_1 , splitterG1ton67n284 , splitterG1ton83n284 , splitterG1ton283n284 , splitterG10ton218n325 , splitterG10ton219n325 , splitterG10ton324n325 , splitterG11ton95n329 , splitterG11ton235n329 , splitterG11ton328n329 , splitterG12ton258n333 , splitterG12ton93n333 , splitterG12ton332n333 , splitterG13ton132n339 , splitterG13ton65n339 , splitterG13ton338n339 , splitterG14ton129n343 , splitterG14ton216n343 , splitterG14ton342n343 , splitterG15ton132n347 , splitterG15ton236n347 , splitterG15ton346n347 , splitterG16ton129n351 , splitterG16ton262n351 , splitterG16ton350n351 , splitterG17ton161n364 , splitterG17ton44n364 , splitterG17ton363n364 , splitterG18ton177n368 , splitterG18ton47n368 , splitterG18ton367n368 , splitterG19ton101n372 , splitterG19ton44n372 , splitterG19ton371n372 , splitterG2ton215n288 , splitterG2ton216n288 , splitterG2ton287n288 , splitterG20ton138n376 , splitterG20ton47n376 , splitterG20ton375n376 , splitterG21ton158n382 , splitterG21ton59n382 , splitterG21ton381n382 , splitterG22ton180n386 , splitterG22ton56n386 , splitterG22ton385n386 , splitterG23ton101n390 , splitterG23ton56n390 , splitterG23ton389n390 , splitterG24ton138n394 , splitterG24ton59n394 , splitterG24ton393n394 , splitterG25ton158n399 , splitterG25ton207n399 , splitterG25ton398n399 , splitterG26ton177n403 , splitterG26ton210n403 , splitterG26ton402n403 , splitterG27ton104n407 , splitterG27ton210n407 , splitterG27ton406n407 , splitterG28ton141n411 , splitterG28ton207n411 , splitterG28ton410n411 , splitterG29ton161n417 , splitterG29ton195n417 , splitterG29ton416n417 , splitterG3ton79n292 , splitterG3ton239n292 , splitterG3ton291n292 , splitterG30ton180n421 , splitterG30ton195n421 , splitterG30ton420n421 , splitterG31ton104n425 , splitterG31ton198n425 , splitterG31ton424n425 , splitterG32ton141n429 , splitterG32ton198n429 , splitterG32ton428n429 , splitterG4ton258n296 , splitterG4ton80n296 , splitterG4ton295n296 , splitterG41ton173n231 , splitterG41ton125n231 , splitterG41ton254n231 , splitterG5ton119n302 , splitterG5ton65n302 , splitterG5ton301n302 , splitterG6ton119n306 , splitterG6ton219n306 , splitterG6ton305n306 , splitterG7ton116n310 , splitterG7ton239n310 , splitterG7ton309n310 , splitterG8ton116n314 , splitterG8ton262n314 , splitterG8ton313n314 , splitterG9ton67n321 , splitterG9ton96n321 , splitterG9ton320n321 , splitterfromn42 , splitterfromn45 , splitterfromn48 , splittern51ton232n53 , splitterfromn54 , splitterfromn57 , splitterfromn60 , splittern63ton255n74 , splitterfromn66 , splitterfromn69 , splitterfromn72 , splitterfromn75 , splittern78ton230n300 , splittern78ton277n300 , splittern78ton337n300 , splittern78ton319n300 , splitterfromn81 , splitterfromn84 , splittern87ton155n90 , splitterfromn88 , splitterfromn91 , splitterfromn94 , splitterfromn97 , splittern100ton110n175 , splitterfromn103 , splitterfromn106 , splitterfromn109 , splitterfromn112 , splittern115ton153n405 , splittern115ton354n405 , splittern115ton388n405 , splittern115ton370n405 , splitterfromn118 , splitterfromn121 , splittern124ton126n168 , splitterfromn125 , splitterfromn128 , splitterfromn131 , splitterfromn134 , splittern137ton147n187 , splitterfromn140 , splitterfromn143 , splitterfromn146 , splitterfromn149 , splittern152ton153n409 , splittern152ton354n409 , splittern152ton392n409 , splittern152ton374n409 , splittern153ton356n281 , splittern153ton317n281 , splitterfromn154 , splitterfromn157 , splitterfromn160 , splitterfromn163 , splitterfromn166 , splitterfromn169 , splittern172ton192n397 , splittern172ton357n397 , splittern172ton380n397 , splittern172ton362n397 , splitterfromn173 , splitterfromn176 , splitterfromn179 , splitterfromn182 , splitterfromn185 , splitterfromn188 , splittern191ton192n401 , splittern191ton357n401 , splittern191ton384n401 , splittern191ton366n401 , splitterfromn192 , splitterfromn193 , splitterfromn196 , splitterfromn199 , splittern202ton203n268 , splitterfromn205 , splitterfromn208 , splitterfromn211 , splittern214ton224n245 , splitterfromn217 , splitterfromn220 , splitterfromn223 , splitterfromn226 , splittern229ton230n304 , splittern229ton277n304 , splittern229ton341n304 , splittern229ton323n304 , splitterfromn230 , splitterfromn231 , splitterfromn234 , splitterfromn237 , splitterfromn240 , splitterfromn243 , splitterfromn246 , splittern249ton250n308 , splittern249ton275n308 , splittern249ton345n308 , splittern249ton327n308 , splitterfromn250 , splitterfromn251 , splitterfromn252 , splitterfromn254 , splitterfromn257 , splitterfromn260 , splitterfromn263 , splitterfromn266 , splitterfromn269 , splittern272ton274n312 , splittern272ton275n312 , splittern272ton273n312 , splittern272ton349n312 , splittern272ton331n312 , splitterfromn274 , splittern279ton280n336 , splitterfromn280 , splittern281ton282n294 , splitterfromn282 , splitterfromn286 , splitterfromn290 , splitterfromn294 , splittern298ton356n299 , splittern298ton335n299 , splittern299ton300n312 , splitterfromn300 , splitterfromn304 , splitterfromn308 , splitterfromn312 , splittern316ton353n318 , splittern316ton335n318 , splittern318ton319n331 , splitterfromn319 , splitterfromn323 , splitterfromn327 , splitterfromn331 , splittern336ton337n349 , splitterfromn337 , splitterfromn341 , splitterfromn345 , splitterfromn349 , splittern359ton360n414 , splitterfromn360 , splittern361ton362n374 , splitterfromn362 , splitterfromn366 , splitterfromn370 , splitterfromn374 , splittern379ton380n392 , splitterfromn380 , splitterfromn384 , splitterfromn388 , splitterfromn392 , splittern396ton397n409 , splitterfromn397 , splitterfromn401 , splitterfromn405 , splitterfromn409 , splittern414ton415n427 , splitterfromn415 , splitterfromn419 , splitterfromn423 , splitterfromn427 ;

PI_AQFP G1_( clk_1 , G1 );
PI_AQFP G10_( clk_1 , G10 );
PI_AQFP G11_( clk_1 , G11 );
PI_AQFP G12_( clk_1 , G12 );
PI_AQFP G13_( clk_1 , G13 );
PI_AQFP G14_( clk_1 , G14 );
PI_AQFP G15_( clk_1 , G15 );
PI_AQFP G16_( clk_1 , G16 );
PI_AQFP G17_( clk_1 , G17 );
PI_AQFP G18_( clk_1 , G18 );
PI_AQFP G19_( clk_1 , G19 );
PI_AQFP G2_( clk_1 , G2 );
PI_AQFP G20_( clk_1 , G20 );
PI_AQFP G21_( clk_1 , G21 );
PI_AQFP G22_( clk_1 , G22 );
PI_AQFP G23_( clk_1 , G23 );
PI_AQFP G24_( clk_1 , G24 );
PI_AQFP G25_( clk_1 , G25 );
PI_AQFP G26_( clk_1 , G26 );
PI_AQFP G27_( clk_1 , G27 );
PI_AQFP G28_( clk_1 , G28 );
PI_AQFP G29_( clk_1 , G29 );
PI_AQFP G3_( clk_1 , G3 );
PI_AQFP G30_( clk_1 , G30 );
PI_AQFP G31_( clk_1 , G31 );
PI_AQFP G32_( clk_1 , G32 );
PI_AQFP G33_( clk_1 , G33 );
PI_AQFP G34_( clk_1 , G34 );
PI_AQFP G35_( clk_1 , G35 );
PI_AQFP G36_( clk_1 , G36 );
PI_AQFP G37_( clk_1 , G37 );
PI_AQFP G38_( clk_1 , G38 );
PI_AQFP G39_( clk_1 , G39 );
PI_AQFP G4_( clk_1 , G4 );
PI_AQFP G40_( clk_1 , G40 );
PI_AQFP G41_( clk_1 , G41 );
PI_AQFP G5_( clk_1 , G5 );
PI_AQFP G6_( clk_1 , G6 );
PI_AQFP G7_( clk_1 , G7 );
PI_AQFP G8_( clk_1 , G8 );
PI_AQFP G9_( clk_1 , G9 );
and_AQFP n42_( clk_5 , buf_G33_n42_1 , splitterG41ton254n231 , 0 , 0 , n42 );
or_AQFP n43_( clk_3 , splitterG17ton161n364 , splitterG19ton101n372 , 0 , 0 , n43 );
and_AQFP n44_( clk_4 , splitterG17ton44n364 , splitterG19ton44n372 , 0 , 0 , n44 );
and_AQFP n45_( clk_5 , n43 , n44 , 0 , 1 , n45 );
and_AQFP n46_( clk_3 , splitterG18ton177n368 , splitterG20ton138n376 , 1 , 0 , n46 );
and_AQFP n47_( clk_4 , splitterG18ton47n368 , splitterG20ton47n376 , 0 , 1 , n47 );
or_AQFP n48_( clk_5 , n46 , n47 , 0 , 0 , n48 );
and_AQFP n49_( clk_7 , splitterfromn45 , splitterfromn48 , 1 , 0 , n49 );
and_AQFP n50_( clk_7 , splitterfromn45 , splitterfromn48 , 0 , 1 , n50 );
or_AQFP n51_( clk_8 , n49 , n50 , 0 , 0 , n51 );
and_AQFP n52_( clk_2 , splitterfromn42 , splittern51ton232n53 , 1 , 0 , n52 );
and_AQFP n53_( clk_2 , splitterfromn42 , splittern51ton232n53 , 0 , 1 , n53 );
or_AQFP n54_( clk_3 , n52 , n53 , 0 , 0 , n54 );
or_AQFP n55_( clk_3 , splitterG22ton180n386 , splitterG23ton101n390 , 0 , 0 , n55 );
and_AQFP n56_( clk_4 , splitterG22ton56n386 , splitterG23ton56n390 , 0 , 0 , n56 );
and_AQFP n57_( clk_5 , n55 , n56 , 0 , 1 , n57 );
and_AQFP n58_( clk_3 , splitterG21ton158n382 , splitterG24ton138n394 , 0 , 1 , n58 );
and_AQFP n59_( clk_4 , splitterG21ton59n382 , splitterG24ton59n394 , 1 , 0 , n59 );
or_AQFP n60_( clk_5 , n58 , n59 , 0 , 0 , n60 );
and_AQFP n61_( clk_7 , splitterfromn57 , splitterfromn60 , 1 , 0 , n61 );
and_AQFP n62_( clk_7 , splitterfromn57 , splitterfromn60 , 0 , 1 , n62 );
or_AQFP n63_( clk_8 , n61 , n62 , 0 , 0 , n63 );
or_AQFP n64_( clk_3 , splitterG13ton132n339 , splitterG5ton119n302 , 0 , 0 , n64 );
and_AQFP n65_( clk_4 , splitterG13ton65n339 , splitterG5ton65n302 , 0 , 0 , n65 );
and_AQFP n66_( clk_5 , n64 , n65 , 0 , 1 , n66 );
and_AQFP n67_( clk_3 , splitterG1ton67n284 , splitterG9ton67n321 , 0 , 1 , n67 );
and_AQFP n68_( clk_3 , splitterG1ton67n284 , splitterG9ton67n321 , 1 , 0 , n68 );
or_AQFP n69_( clk_4 , n67 , n68 , 0 , 0 , n69 );
or_AQFP n70_( clk_7 , splitterfromn66 , splitterfromn69 , 0 , 0 , n70 );
and_AQFP n71_( clk_7 , splitterfromn66 , splitterfromn69 , 0 , 0 , n71 );
and_AQFP n72_( clk_8 , n70 , n71 , 0 , 1 , n72 );
and_AQFP n73_( clk_2 , splittern63ton255n74 , splitterfromn72 , 0 , 0 , n73 );
or_AQFP n74_( clk_2 , splittern63ton255n74 , splitterfromn72 , 0 , 0 , n74 );
and_AQFP n75_( clk_3 , n73 , n74 , 1 , 0 , n75 );
and_AQFP n76_( clk_5 , splitterfromn54 , splitterfromn75 , 1 , 0 , n76 );
and_AQFP n77_( clk_5 , splitterfromn54 , splitterfromn75 , 0 , 1 , n77 );
or_AQFP n78_( clk_6 , n76 , n77 , 0 , 0 , n78 );
or_AQFP n79_( clk_3 , splitterG3ton79n292 , splitterG4ton258n296 , 0 , 0 , n79 );
and_AQFP n80_( clk_4 , splitterG3ton79n292 , splitterG4ton80n296 , 0 , 0 , n80 );
and_AQFP n81_( clk_5 , n79 , n80 , 0 , 1 , n81 );
and_AQFP n82_( clk_3 , splitterG1ton67n284 , splitterG2ton215n288 , 0 , 1 , n82 );
and_AQFP n83_( clk_4 , splitterG1ton83n284 , splitterG2ton216n288 , 1 , 0 , n83 );
or_AQFP n84_( clk_5 , n82 , n83 , 0 , 0 , n84 );
and_AQFP n85_( clk_7 , splitterfromn81 , splitterfromn84 , 1 , 0 , n85 );
and_AQFP n86_( clk_7 , splitterfromn81 , splitterfromn84 , 0 , 1 , n86 );
or_AQFP n87_( clk_8 , n85 , n86 , 0 , 0 , n87 );
and_AQFP n88_( clk_5 , buf_G39_n88_1 , splitterG41ton254n231 , 0 , 0 , n88 );
and_AQFP n89_( clk_2 , splittern87ton155n90 , splitterfromn88 , 0 , 1 , n89 );
and_AQFP n90_( clk_2 , splittern87ton155n90 , splitterfromn88 , 1 , 0 , n90 );
or_AQFP n91_( clk_3 , n89 , n90 , 0 , 0 , n91 );
or_AQFP n92_( clk_3 , splitterG10ton218n325 , splitterG12ton258n333 , 0 , 0 , n92 );
and_AQFP n93_( clk_4 , splitterG10ton219n325 , splitterG12ton93n333 , 0 , 0 , n93 );
and_AQFP n94_( clk_5 , n92 , n93 , 0 , 1 , n94 );
and_AQFP n95_( clk_3 , splitterG11ton95n329 , splitterG9ton67n321 , 1 , 0 , n95 );
and_AQFP n96_( clk_4 , splitterG11ton235n329 , splitterG9ton96n321 , 0 , 1 , n96 );
or_AQFP n97_( clk_5 , n95 , n96 , 0 , 0 , n97 );
and_AQFP n98_( clk_7 , splitterfromn94 , splitterfromn97 , 1 , 0 , n98 );
and_AQFP n99_( clk_7 , splitterfromn94 , splitterfromn97 , 0 , 1 , n99 );
or_AQFP n100_( clk_8 , n98 , n99 , 0 , 0 , n100 );
or_AQFP n101_( clk_3 , splitterG19ton101n372 , splitterG23ton101n390 , 0 , 0 , n101 );
and_AQFP n102_( clk_3 , splitterG19ton101n372 , splitterG23ton101n390 , 0 , 0 , n102 );
and_AQFP n103_( clk_4 , n101 , n102 , 0 , 1 , n103 );
and_AQFP n104_( clk_3 , splitterG27ton104n407 , splitterG31ton104n425 , 0 , 1 , n104 );
and_AQFP n105_( clk_3 , splitterG27ton104n407 , splitterG31ton104n425 , 1 , 0 , n105 );
or_AQFP n106_( clk_4 , n104 , n105 , 0 , 0 , n106 );
or_AQFP n107_( clk_6 , splitterfromn103 , splitterfromn106 , 0 , 0 , n107 );
and_AQFP n108_( clk_6 , splitterfromn103 , splitterfromn106 , 0 , 0 , n108 );
and_AQFP n109_( clk_7 , n107 , n108 , 0 , 1 , n109 );
and_AQFP n110_( clk_2 , splittern100ton110n175 , splitterfromn109 , 0 , 0 , n110 );
or_AQFP n111_( clk_2 , splittern100ton110n175 , splitterfromn109 , 0 , 0 , n111 );
and_AQFP n112_( clk_3 , n110 , n111 , 1 , 0 , n112 );
and_AQFP n113_( clk_5 , splitterfromn91 , splitterfromn112 , 1 , 0 , n113 );
and_AQFP n114_( clk_5 , splitterfromn91 , splitterfromn112 , 0 , 1 , n114 );
or_AQFP n115_( clk_6 , n113 , n114 , 0 , 0 , n115 );
or_AQFP n116_( clk_3 , splitterG7ton116n310 , splitterG8ton116n314 , 0 , 0 , n116 );
and_AQFP n117_( clk_3 , splitterG7ton116n310 , splitterG8ton116n314 , 0 , 0 , n117 );
and_AQFP n118_( clk_4 , n116 , n117 , 0 , 1 , n118 );
and_AQFP n119_( clk_3 , splitterG5ton119n302 , splitterG6ton119n306 , 1 , 0 , n119 );
and_AQFP n120_( clk_3 , splitterG5ton119n302 , splitterG6ton119n306 , 0 , 1 , n120 );
or_AQFP n121_( clk_4 , n119 , n120 , 0 , 0 , n121 );
and_AQFP n122_( clk_6 , splitterfromn118 , splitterfromn121 , 1 , 0 , n122 );
and_AQFP n123_( clk_6 , splitterfromn118 , splitterfromn121 , 0 , 1 , n123 );
or_AQFP n124_( clk_7 , n122 , n123 , 0 , 0 , n124 );
and_AQFP n125_( clk_4 , buf_G40_n125_1 , splitterG41ton125n231 , 0 , 0 , n125 );
and_AQFP n126_( clk_1 , splittern124ton126n168 , splitterfromn125 , 0 , 1 , n126 );
and_AQFP n127_( clk_1 , splittern124ton126n168 , splitterfromn125 , 1 , 0 , n127 );
or_AQFP n128_( clk_2 , n126 , n127 , 0 , 0 , n128 );
or_AQFP n129_( clk_3 , splitterG14ton129n343 , splitterG16ton129n351 , 0 , 0 , n129 );
and_AQFP n130_( clk_3 , splitterG14ton129n343 , splitterG16ton129n351 , 0 , 0 , n130 );
and_AQFP n131_( clk_4 , n129 , n130 , 0 , 1 , n131 );
and_AQFP n132_( clk_3 , splitterG13ton132n339 , splitterG15ton132n347 , 0 , 1 , n132 );
and_AQFP n133_( clk_3 , splitterG13ton132n339 , splitterG15ton132n347 , 1 , 0 , n133 );
or_AQFP n134_( clk_4 , n132 , n133 , 0 , 0 , n134 );
and_AQFP n135_( clk_6 , splitterfromn131 , splitterfromn134 , 1 , 0 , n135 );
and_AQFP n136_( clk_6 , splitterfromn131 , splitterfromn134 , 0 , 1 , n136 );
or_AQFP n137_( clk_7 , n135 , n136 , 0 , 0 , n137 );
or_AQFP n138_( clk_3 , splitterG20ton138n376 , splitterG24ton138n394 , 0 , 0 , n138 );
and_AQFP n139_( clk_3 , splitterG20ton138n376 , splitterG24ton138n394 , 0 , 0 , n139 );
and_AQFP n140_( clk_4 , n138 , n139 , 0 , 1 , n140 );
and_AQFP n141_( clk_3 , splitterG28ton141n411 , splitterG32ton141n429 , 1 , 0 , n141 );
and_AQFP n142_( clk_3 , splitterG28ton141n411 , splitterG32ton141n429 , 0 , 1 , n142 );
or_AQFP n143_( clk_4 , n141 , n142 , 0 , 0 , n143 );
or_AQFP n144_( clk_6 , splitterfromn140 , splitterfromn143 , 0 , 0 , n144 );
and_AQFP n145_( clk_6 , splitterfromn140 , splitterfromn143 , 0 , 0 , n145 );
and_AQFP n146_( clk_7 , n144 , n145 , 0 , 1 , n146 );
and_AQFP n147_( clk_1 , splittern137ton147n187 , splitterfromn146 , 0 , 0 , n147 );
or_AQFP n148_( clk_1 , splittern137ton147n187 , splitterfromn146 , 0 , 0 , n148 );
and_AQFP n149_( clk_2 , n147 , n148 , 1 , 0 , n149 );
and_AQFP n150_( clk_5 , splitterfromn128 , splitterfromn149 , 1 , 0 , n150 );
and_AQFP n151_( clk_5 , splitterfromn128 , splitterfromn149 , 0 , 1 , n151 );
or_AQFP n152_( clk_6 , n150 , n151 , 0 , 0 , n152 );
and_AQFP n153_( clk_8 , splittern115ton153n405 , splittern152ton153n409 , 0 , 1 , n153 );
and_AQFP n154_( clk_4 , buf_G37_n154_1 , splitterG41ton125n231 , 0 , 0 , n154 );
and_AQFP n155_( clk_2 , splittern87ton155n90 , splitterfromn154 , 0 , 1 , n155 );
and_AQFP n156_( clk_2 , splittern87ton155n90 , splitterfromn154 , 1 , 0 , n156 );
or_AQFP n157_( clk_3 , n155 , n156 , 0 , 0 , n157 );
and_AQFP n158_( clk_3 , splitterG21ton158n382 , splitterG25ton158n399 , 0 , 1 , n158 );
and_AQFP n159_( clk_3 , splitterG21ton158n382 , splitterG25ton158n399 , 1 , 0 , n159 );
or_AQFP n160_( clk_4 , n158 , n159 , 0 , 0 , n160 );
or_AQFP n161_( clk_3 , splitterG17ton161n364 , splitterG29ton161n417 , 0 , 0 , n161 );
and_AQFP n162_( clk_3 , splitterG17ton161n364 , splitterG29ton161n417 , 0 , 0 , n162 );
and_AQFP n163_( clk_4 , n161 , n162 , 0 , 1 , n163 );
or_AQFP n164_( clk_6 , splitterfromn160 , splitterfromn163 , 0 , 0 , n164 );
and_AQFP n165_( clk_6 , splitterfromn160 , splitterfromn163 , 0 , 0 , n165 );
and_AQFP n166_( clk_7 , n164 , n165 , 0 , 1 , n166 );
and_AQFP n167_( clk_1 , splittern124ton126n168 , splitterfromn166 , 0 , 0 , n167 );
or_AQFP n168_( clk_1 , splittern124ton126n168 , splitterfromn166 , 0 , 0 , n168 );
and_AQFP n169_( clk_3 , n167 , n168 , 1 , 0 , n169 );
and_AQFP n170_( clk_5 , splitterfromn157 , splitterfromn169 , 1 , 0 , n170 );
and_AQFP n171_( clk_5 , splitterfromn157 , splitterfromn169 , 0 , 1 , n171 );
or_AQFP n172_( clk_6 , n170 , n171 , 0 , 0 , n172 );
and_AQFP n173_( clk_3 , G38 , splitterG41ton173n231 , 0 , 0 , n173 );
and_AQFP n174_( clk_2 , splittern100ton110n175 , splitterfromn173 , 0 , 1 , n174 );
and_AQFP n175_( clk_2 , splittern100ton110n175 , splitterfromn173 , 1 , 0 , n175 );
or_AQFP n176_( clk_3 , n174 , n175 , 0 , 0 , n176 );
and_AQFP n177_( clk_3 , splitterG18ton177n368 , splitterG26ton177n403 , 1 , 0 , n177 );
and_AQFP n178_( clk_3 , splitterG18ton177n368 , splitterG26ton177n403 , 0 , 1 , n178 );
or_AQFP n179_( clk_4 , n177 , n178 , 0 , 0 , n179 );
or_AQFP n180_( clk_3 , splitterG22ton180n386 , splitterG30ton180n421 , 0 , 0 , n180 );
and_AQFP n181_( clk_3 , splitterG22ton180n386 , splitterG30ton180n421 , 0 , 0 , n181 );
and_AQFP n182_( clk_4 , n180 , n181 , 0 , 1 , n182 );
or_AQFP n183_( clk_6 , splitterfromn179 , splitterfromn182 , 0 , 0 , n183 );
and_AQFP n184_( clk_6 , splitterfromn179 , splitterfromn182 , 0 , 0 , n184 );
and_AQFP n185_( clk_7 , n183 , n184 , 0 , 1 , n185 );
and_AQFP n186_( clk_1 , splittern137ton147n187 , splitterfromn185 , 0 , 0 , n186 );
or_AQFP n187_( clk_1 , splittern137ton147n187 , splitterfromn185 , 0 , 0 , n187 );
and_AQFP n188_( clk_2 , n186 , n187 , 1 , 0 , n188 );
and_AQFP n189_( clk_5 , splitterfromn176 , splitterfromn188 , 1 , 0 , n189 );
and_AQFP n190_( clk_5 , splitterfromn176 , splitterfromn188 , 0 , 1 , n190 );
or_AQFP n191_( clk_6 , n189 , n190 , 0 , 0 , n191 );
and_AQFP n192_( clk_8 , splittern172ton192n397 , splittern191ton192n401 , 0 , 1 , n192 );
and_AQFP n193_( clk_4 , buf_G34_n193_1 , splitterG41ton125n231 , 0 , 0 , n193 );
or_AQFP n194_( clk_3 , splitterG29ton161n417 , splitterG30ton180n421 , 0 , 0 , n194 );
and_AQFP n195_( clk_4 , splitterG29ton195n417 , splitterG30ton195n421 , 0 , 0 , n195 );
and_AQFP n196_( clk_5 , n194 , n195 , 0 , 1 , n196 );
and_AQFP n197_( clk_3 , splitterG31ton104n425 , splitterG32ton141n429 , 1 , 0 , n197 );
and_AQFP n198_( clk_4 , splitterG31ton198n425 , splitterG32ton198n429 , 0 , 1 , n198 );
or_AQFP n199_( clk_5 , n197 , n198 , 0 , 0 , n199 );
and_AQFP n200_( clk_7 , splitterfromn196 , splitterfromn199 , 1 , 0 , n200 );
and_AQFP n201_( clk_7 , splitterfromn196 , splitterfromn199 , 0 , 1 , n201 );
or_AQFP n202_( clk_8 , n200 , n201 , 0 , 0 , n202 );
and_AQFP n203_( clk_2 , splitterfromn193 , splittern202ton203n268 , 1 , 0 , n203 );
and_AQFP n204_( clk_2 , splitterfromn193 , splittern202ton203n268 , 0 , 1 , n204 );
or_AQFP n205_( clk_3 , n203 , n204 , 0 , 0 , n205 );
or_AQFP n206_( clk_3 , splitterG25ton158n399 , splitterG28ton141n411 , 0 , 0 , n206 );
and_AQFP n207_( clk_4 , splitterG25ton207n399 , splitterG28ton207n411 , 0 , 0 , n207 );
and_AQFP n208_( clk_5 , n206 , n207 , 0 , 1 , n208 );
and_AQFP n209_( clk_3 , splitterG26ton177n403 , splitterG27ton104n407 , 0 , 1 , n209 );
and_AQFP n210_( clk_4 , splitterG26ton210n403 , splitterG27ton210n407 , 1 , 0 , n210 );
or_AQFP n211_( clk_5 , n209 , n210 , 0 , 0 , n211 );
and_AQFP n212_( clk_7 , splitterfromn208 , splitterfromn211 , 1 , 0 , n212 );
and_AQFP n213_( clk_7 , splitterfromn208 , splitterfromn211 , 0 , 1 , n213 );
or_AQFP n214_( clk_8 , n212 , n213 , 0 , 0 , n214 );
or_AQFP n215_( clk_3 , splitterG14ton129n343 , splitterG2ton215n288 , 0 , 0 , n215 );
and_AQFP n216_( clk_4 , splitterG14ton216n343 , splitterG2ton216n288 , 0 , 0 , n216 );
and_AQFP n217_( clk_5 , n215 , n216 , 0 , 1 , n217 );
and_AQFP n218_( clk_3 , splitterG10ton218n325 , splitterG6ton119n306 , 0 , 1 , n218 );
and_AQFP n219_( clk_4 , splitterG10ton219n325 , splitterG6ton219n306 , 1 , 0 , n219 );
or_AQFP n220_( clk_5 , n218 , n219 , 0 , 0 , n220 );
or_AQFP n221_( clk_7 , splitterfromn217 , splitterfromn220 , 0 , 0 , n221 );
and_AQFP n222_( clk_7 , splitterfromn217 , splitterfromn220 , 0 , 0 , n222 );
and_AQFP n223_( clk_8 , n221 , n222 , 0 , 1 , n223 );
and_AQFP n224_( clk_2 , splittern214ton224n245 , splitterfromn223 , 0 , 0 , n224 );
or_AQFP n225_( clk_2 , splittern214ton224n245 , splitterfromn223 , 0 , 0 , n225 );
and_AQFP n226_( clk_3 , n224 , n225 , 1 , 0 , n226 );
and_AQFP n227_( clk_5 , splitterfromn205 , splitterfromn226 , 1 , 0 , n227 );
and_AQFP n228_( clk_5 , splitterfromn205 , splitterfromn226 , 0 , 1 , n228 );
or_AQFP n229_( clk_6 , n227 , n228 , 0 , 0 , n229 );
and_AQFP n230_( clk_8 , splittern78ton230n300 , splittern229ton230n304 , 1 , 0 , n230 );
and_AQFP n231_( clk_5 , buf_G35_n231_1 , splitterG41ton254n231 , 0 , 0 , n231 );
and_AQFP n232_( clk_2 , splittern51ton232n53 , splitterfromn231 , 0 , 1 , n232 );
and_AQFP n233_( clk_2 , splittern51ton232n53 , splitterfromn231 , 1 , 0 , n233 );
or_AQFP n234_( clk_3 , n232 , n233 , 0 , 0 , n234 );
and_AQFP n235_( clk_4 , splitterG11ton235n329 , splitterG15ton132n347 , 0 , 1 , n235 );
and_AQFP n236_( clk_5 , splitterG11ton235n329 , splitterG15ton236n347 , 1 , 0 , n236 );
or_AQFP n237_( clk_6 , n235 , n236 , 0 , 0 , n237 );
or_AQFP n238_( clk_4 , splitterG3ton79n292 , splitterG7ton116n310 , 0 , 0 , n238 );
and_AQFP n239_( clk_5 , splitterG3ton239n292 , splitterG7ton239n310 , 0 , 0 , n239 );
and_AQFP n240_( clk_6 , n238 , n239 , 0 , 1 , n240 );
or_AQFP n241_( clk_8 , splitterfromn237 , splitterfromn240 , 0 , 0 , n241 );
and_AQFP n242_( clk_8 , splitterfromn237 , splitterfromn240 , 0 , 0 , n242 );
and_AQFP n243_( clk_1 , n241 , n242 , 0 , 1 , n243 );
and_AQFP n244_( clk_3 , splittern214ton224n245 , splitterfromn243 , 0 , 0 , n244 );
or_AQFP n245_( clk_3 , splittern214ton224n245 , splitterfromn243 , 0 , 0 , n245 );
and_AQFP n246_( clk_4 , n244 , n245 , 1 , 0 , n246 );
and_AQFP n247_( clk_6 , splitterfromn234 , splitterfromn246 , 1 , 0 , n247 );
and_AQFP n248_( clk_6 , splitterfromn234 , splitterfromn246 , 0 , 1 , n248 );
or_AQFP n249_( clk_7 , n247 , n248 , 0 , 0 , n249 );
and_AQFP n250_( clk_2 , splitterfromn230 , splittern249ton250n308 , 0 , 1 , n250 );
and_AQFP n251_( clk_8 , splittern78ton230n300 , splittern229ton230n304 , 0 , 1 , n251 );
and_AQFP n252_( clk_2 , splittern249ton250n308 , splitterfromn251 , 1 , 0 , n252 );
or_AQFP n253_( clk_4 , splitterfromn250 , splitterfromn252 , 0 , 0 , n253 );
and_AQFP n254_( clk_5 , buf_G36_n254_1 , splitterG41ton254n231 , 0 , 0 , n254 );
and_AQFP n255_( clk_2 , splittern63ton255n74 , splitterfromn254 , 0 , 1 , n255 );
and_AQFP n256_( clk_2 , splittern63ton255n74 , splitterfromn254 , 1 , 0 , n256 );
or_AQFP n257_( clk_3 , n255 , n256 , 0 , 0 , n257 );
and_AQFP n258_( clk_3 , splitterG12ton258n333 , splitterG4ton258n296 , 0 , 1 , n258 );
and_AQFP n259_( clk_3 , splitterG12ton258n333 , splitterG4ton258n296 , 1 , 0 , n259 );
or_AQFP n260_( clk_4 , n258 , n259 , 0 , 0 , n260 );
or_AQFP n261_( clk_4 , splitterG16ton129n351 , splitterG8ton116n314 , 0 , 0 , n261 );
and_AQFP n262_( clk_5 , splitterG16ton262n351 , splitterG8ton262n314 , 0 , 0 , n262 );
and_AQFP n263_( clk_6 , n261 , n262 , 0 , 1 , n263 );
or_AQFP n264_( clk_8 , splitterfromn260 , splitterfromn263 , 0 , 0 , n264 );
and_AQFP n265_( clk_8 , splitterfromn260 , splitterfromn263 , 0 , 0 , n265 );
and_AQFP n266_( clk_1 , n264 , n265 , 0 , 1 , n266 );
and_AQFP n267_( clk_3 , splittern202ton203n268 , splitterfromn266 , 0 , 0 , n267 );
or_AQFP n268_( clk_3 , splittern202ton203n268 , splitterfromn266 , 0 , 0 , n268 );
and_AQFP n269_( clk_4 , n267 , n268 , 1 , 0 , n269 );
and_AQFP n270_( clk_6 , splitterfromn257 , splitterfromn269 , 1 , 0 , n270 );
and_AQFP n271_( clk_6 , splitterfromn257 , splitterfromn269 , 0 , 1 , n271 );
or_AQFP n272_( clk_7 , n270 , n271 , 0 , 0 , n272 );
and_AQFP n273_( clk_5 , n253 , splittern272ton273n312 , 0 , 1 , n273 );
and_AQFP n274_( clk_2 , splittern249ton250n308 , splittern272ton274n312 , 0 , 1 , n274 );
and_AQFP n275_( clk_3 , splittern249ton275n308 , splittern272ton275n312 , 1 , 0 , n275 );
or_AQFP n276_( clk_4 , splitterfromn274 , n275 , 0 , 0 , n276 );
or_AQFP n277_( clk_3 , splittern78ton277n300 , splittern229ton277n304 , 0 , 0 , n277 );
and_AQFP n278_( clk_5 , n276 , n277 , 0 , 1 , n278 );
or_AQFP n279_( clk_6 , n273 , n278 , 0 , 0 , n279 );
and_AQFP n280_( clk_8 , buf_splitterfromn192_n280_1 , splittern279ton280n336 , 0 , 0 , n280 );
and_AQFP n281_( clk_2 , buf_splittern153ton317n281_n281_1 , splitterfromn280 , 0 , 0 , n281 );
and_AQFP n282_( clk_4 , splittern78ton319n300 , splittern281ton282n294 , 0 , 0 , n282 );
and_AQFP n283_( clk_6 , splitterG1ton283n284 , splitterfromn282 , 0 , 1 , n283 );
and_AQFP n284_( clk_6 , splitterG1ton283n284 , splitterfromn282 , 1 , 0 , n284 );
or_AQFP n285_( clk_7 , n283 , n284 , 0 , 0 , n285 );
and_AQFP n286_( clk_4 , splittern229ton323n304 , splittern281ton282n294 , 0 , 0 , n286 );
and_AQFP n287_( clk_6 , splitterG2ton287n288 , splitterfromn286 , 0 , 1 , n287 );
and_AQFP n288_( clk_6 , splitterG2ton287n288 , splitterfromn286 , 1 , 0 , n288 );
or_AQFP n289_( clk_7 , n287 , n288 , 0 , 0 , n289 );
and_AQFP n290_( clk_4 , splittern249ton327n308 , splittern281ton282n294 , 0 , 0 , n290 );
and_AQFP n291_( clk_6 , splitterG3ton291n292 , splitterfromn290 , 0 , 1 , n291 );
and_AQFP n292_( clk_6 , splitterG3ton291n292 , splitterfromn290 , 1 , 0 , n292 );
or_AQFP n293_( clk_7 , n291 , n292 , 0 , 0 , n293 );
and_AQFP n294_( clk_4 , splittern272ton331n312 , splittern281ton282n294 , 0 , 0 , n294 );
and_AQFP n295_( clk_6 , splitterG4ton295n296 , splitterfromn294 , 0 , 1 , n295 );
and_AQFP n296_( clk_6 , splitterG4ton295n296 , splitterfromn294 , 1 , 0 , n296 );
or_AQFP n297_( clk_7 , n295 , n296 , 0 , 0 , n297 );
and_AQFP n298_( clk_8 , splittern115ton153n405 , splittern152ton153n409 , 1 , 0 , n298 );
and_AQFP n299_( clk_2 , splitterfromn280 , buf_splittern298ton335n299_n299_1 , 0 , 0 , n299 );
and_AQFP n300_( clk_4 , splittern78ton319n300 , splittern299ton300n312 , 0 , 0 , n300 );
and_AQFP n301_( clk_6 , splitterG5ton301n302 , splitterfromn300 , 0 , 1 , n301 );
and_AQFP n302_( clk_6 , splitterG5ton301n302 , splitterfromn300 , 1 , 0 , n302 );
or_AQFP n303_( clk_7 , n301 , n302 , 0 , 0 , n303 );
and_AQFP n304_( clk_4 , splittern229ton323n304 , splittern299ton300n312 , 0 , 0 , n304 );
and_AQFP n305_( clk_6 , splitterG6ton305n306 , splitterfromn304 , 0 , 1 , n305 );
and_AQFP n306_( clk_6 , splitterG6ton305n306 , splitterfromn304 , 1 , 0 , n306 );
or_AQFP n307_( clk_7 , n305 , n306 , 0 , 0 , n307 );
and_AQFP n308_( clk_4 , splittern249ton327n308 , splittern299ton300n312 , 0 , 0 , n308 );
and_AQFP n309_( clk_6 , splitterG7ton309n310 , splitterfromn308 , 0 , 1 , n309 );
and_AQFP n310_( clk_6 , splitterG7ton309n310 , splitterfromn308 , 1 , 0 , n310 );
or_AQFP n311_( clk_7 , n309 , n310 , 0 , 0 , n311 );
and_AQFP n312_( clk_4 , splittern272ton331n312 , splittern299ton300n312 , 0 , 0 , n312 );
and_AQFP n313_( clk_6 , splitterG8ton313n314 , splitterfromn312 , 0 , 1 , n313 );
and_AQFP n314_( clk_6 , splitterG8ton313n314 , splitterfromn312 , 1 , 0 , n314 );
or_AQFP n315_( clk_7 , n313 , n314 , 0 , 0 , n315 );
and_AQFP n316_( clk_8 , splittern172ton192n397 , splittern191ton192n401 , 1 , 0 , n316 );
and_AQFP n317_( clk_8 , splittern153ton317n281 , splittern279ton280n336 , 0 , 0 , n317 );
and_AQFP n318_( clk_1 , buf_splittern316ton335n318_n318_1 , n317 , 0 , 0 , n318 );
and_AQFP n319_( clk_3 , splittern78ton319n300 , splittern318ton319n331 , 0 , 0 , n319 );
and_AQFP n320_( clk_5 , splitterG9ton320n321 , splitterfromn319 , 0 , 1 , n320 );
and_AQFP n321_( clk_5 , splitterG9ton320n321 , splitterfromn319 , 1 , 0 , n321 );
or_AQFP n322_( clk_6 , n320 , n321 , 0 , 0 , n322 );
and_AQFP n323_( clk_3 , splittern229ton323n304 , splittern318ton319n331 , 0 , 0 , n323 );
and_AQFP n324_( clk_5 , splitterG10ton324n325 , splitterfromn323 , 0 , 1 , n324 );
and_AQFP n325_( clk_5 , splitterG10ton324n325 , splitterfromn323 , 1 , 0 , n325 );
or_AQFP n326_( clk_6 , n324 , n325 , 0 , 0 , n326 );
and_AQFP n327_( clk_3 , splittern249ton327n308 , splittern318ton319n331 , 0 , 0 , n327 );
and_AQFP n328_( clk_5 , splitterG11ton328n329 , splitterfromn327 , 0 , 1 , n328 );
and_AQFP n329_( clk_5 , splitterG11ton328n329 , splitterfromn327 , 1 , 0 , n329 );
or_AQFP n330_( clk_6 , n328 , n329 , 0 , 0 , n330 );
and_AQFP n331_( clk_3 , splittern272ton331n312 , splittern318ton319n331 , 0 , 0 , n331 );
and_AQFP n332_( clk_5 , splitterG12ton332n333 , splitterfromn331 , 0 , 1 , n332 );
and_AQFP n333_( clk_5 , splitterG12ton332n333 , splitterfromn331 , 1 , 0 , n333 );
or_AQFP n334_( clk_7 , n332 , n333 , 0 , 0 , n334 );
and_AQFP n335_( clk_6 , splittern298ton335n299 , splittern316ton335n318 , 0 , 0 , n335 );
and_AQFP n336_( clk_8 , splittern279ton280n336 , n335 , 0 , 0 , n336 );
and_AQFP n337_( clk_2 , splittern78ton337n300 , splittern336ton337n349 , 0 , 0 , n337 );
or_AQFP n338_( clk_4 , splitterG13ton338n339 , splitterfromn337 , 0 , 0 , n338 );
and_AQFP n339_( clk_4 , splitterG13ton338n339 , splitterfromn337 , 0 , 0 , n339 );
and_AQFP n340_( clk_6 , n338 , n339 , 0 , 1 , n340 );
and_AQFP n341_( clk_2 , splittern229ton341n304 , splittern336ton337n349 , 0 , 0 , n341 );
or_AQFP n342_( clk_4 , splitterG14ton342n343 , splitterfromn341 , 0 , 0 , n342 );
and_AQFP n343_( clk_4 , splitterG14ton342n343 , splitterfromn341 , 0 , 0 , n343 );
and_AQFP n344_( clk_6 , n342 , n343 , 0 , 1 , n344 );
and_AQFP n345_( clk_2 , splittern249ton345n308 , splittern336ton337n349 , 0 , 0 , n345 );
and_AQFP n346_( clk_4 , splitterG15ton346n347 , splitterfromn345 , 0 , 1 , n346 );
and_AQFP n347_( clk_4 , splitterG15ton346n347 , splitterfromn345 , 1 , 0 , n347 );
or_AQFP n348_( clk_6 , n346 , n347 , 0 , 0 , n348 );
and_AQFP n349_( clk_2 , splittern272ton349n312 , splittern336ton337n349 , 0 , 0 , n349 );
or_AQFP n350_( clk_4 , splitterG16ton350n351 , splitterfromn349 , 0 , 0 , n350 );
and_AQFP n351_( clk_4 , splitterG16ton350n351 , splitterfromn349 , 0 , 0 , n351 );
and_AQFP n352_( clk_6 , n350 , n351 , 0 , 1 , n352 );
or_AQFP n353_( clk_2 , splitterfromn192 , splittern316ton353n318 , 0 , 0 , n353 );
or_AQFP n354_( clk_2 , splittern115ton354n405 , splittern152ton354n409 , 0 , 0 , n354 );
and_AQFP n355_( clk_3 , n353 , n354 , 0 , 1 , n355 );
or_AQFP n356_( clk_2 , splittern153ton356n281 , splittern298ton356n299 , 0 , 0 , n356 );
or_AQFP n357_( clk_2 , splittern172ton357n397 , splittern191ton357n401 , 0 , 0 , n357 );
and_AQFP n358_( clk_3 , n356 , n357 , 0 , 1 , n358 );
or_AQFP n359_( clk_4 , n355 , n358 , 0 , 0 , n359 );
and_AQFP n360_( clk_6 , buf_splitterfromn274_n360_1 , splittern359ton360n414 , 0 , 0 , n360 );
and_AQFP n361_( clk_8 , buf_splitterfromn251_n361_1 , splitterfromn360 , 0 , 0 , n361 );
and_AQFP n362_( clk_2 , splittern172ton362n397 , splittern361ton362n374 , 0 , 0 , n362 );
and_AQFP n363_( clk_4 , splitterG17ton363n364 , splitterfromn362 , 0 , 1 , n363 );
and_AQFP n364_( clk_4 , splitterG17ton363n364 , splitterfromn362 , 1 , 0 , n364 );
or_AQFP n365_( clk_6 , n363 , n364 , 0 , 0 , n365 );
and_AQFP n366_( clk_2 , splittern191ton366n401 , splittern361ton362n374 , 0 , 0 , n366 );
and_AQFP n367_( clk_4 , splitterG18ton367n368 , splitterfromn366 , 0 , 1 , n367 );
and_AQFP n368_( clk_4 , splitterG18ton367n368 , splitterfromn366 , 1 , 0 , n368 );
or_AQFP n369_( clk_6 , n367 , n368 , 0 , 0 , n369 );
and_AQFP n370_( clk_2 , splittern115ton370n405 , splittern361ton362n374 , 0 , 0 , n370 );
and_AQFP n371_( clk_4 , splitterG19ton371n372 , splitterfromn370 , 0 , 1 , n371 );
and_AQFP n372_( clk_4 , splitterG19ton371n372 , splitterfromn370 , 1 , 0 , n372 );
or_AQFP n373_( clk_6 , n371 , n372 , 0 , 0 , n373 );
and_AQFP n374_( clk_2 , splittern152ton374n409 , splittern361ton362n374 , 0 , 0 , n374 );
and_AQFP n375_( clk_4 , splitterG20ton375n376 , splitterfromn374 , 0 , 1 , n375 );
and_AQFP n376_( clk_4 , splitterG20ton375n376 , splitterfromn374 , 1 , 0 , n376 );
or_AQFP n377_( clk_6 , n375 , n376 , 0 , 0 , n377 );
and_AQFP n378_( clk_5 , splitterfromn252 , splittern272ton273n312 , 0 , 0 , n378 );
and_AQFP n379_( clk_6 , splittern359ton360n414 , n378 , 0 , 0 , n379 );
and_AQFP n380_( clk_8 , splittern172ton380n397 , splittern379ton380n392 , 0 , 0 , n380 );
and_AQFP n381_( clk_2 , splitterG21ton381n382 , splitterfromn380 , 0 , 1 , n381 );
and_AQFP n382_( clk_2 , splitterG21ton381n382 , splitterfromn380 , 1 , 0 , n382 );
or_AQFP n383_( clk_4 , n381 , n382 , 0 , 0 , n383 );
and_AQFP n384_( clk_8 , splittern191ton384n401 , splittern379ton380n392 , 0 , 0 , n384 );
and_AQFP n385_( clk_2 , splitterG22ton385n386 , splitterfromn384 , 0 , 1 , n385 );
and_AQFP n386_( clk_2 , splitterG22ton385n386 , splitterfromn384 , 1 , 0 , n386 );
or_AQFP n387_( clk_4 , n385 , n386 , 0 , 0 , n387 );
and_AQFP n388_( clk_8 , splittern115ton388n405 , splittern379ton380n392 , 0 , 0 , n388 );
and_AQFP n389_( clk_2 , splitterG23ton389n390 , splitterfromn388 , 0 , 1 , n389 );
and_AQFP n390_( clk_2 , splitterG23ton389n390 , splitterfromn388 , 1 , 0 , n390 );
or_AQFP n391_( clk_4 , n389 , n390 , 0 , 0 , n391 );
and_AQFP n392_( clk_8 , splittern152ton392n409 , splittern379ton380n392 , 0 , 0 , n392 );
and_AQFP n393_( clk_2 , splitterG24ton393n394 , splitterfromn392 , 0 , 1 , n393 );
and_AQFP n394_( clk_2 , splitterG24ton393n394 , splitterfromn392 , 1 , 0 , n394 );
or_AQFP n395_( clk_4 , n393 , n394 , 0 , 0 , n395 );
and_AQFP n396_( clk_8 , buf_splitterfromn230_n396_1 , splitterfromn360 , 0 , 0 , n396 );
and_AQFP n397_( clk_2 , splittern172ton362n397 , splittern396ton397n409 , 0 , 0 , n397 );
and_AQFP n398_( clk_4 , splitterG25ton398n399 , splitterfromn397 , 0 , 1 , n398 );
and_AQFP n399_( clk_4 , splitterG25ton398n399 , splitterfromn397 , 1 , 0 , n399 );
or_AQFP n400_( clk_6 , n398 , n399 , 0 , 0 , n400 );
and_AQFP n401_( clk_2 , splittern191ton366n401 , splittern396ton397n409 , 0 , 0 , n401 );
and_AQFP n402_( clk_4 , splitterG26ton402n403 , splitterfromn401 , 0 , 1 , n402 );
and_AQFP n403_( clk_4 , splitterG26ton402n403 , splitterfromn401 , 1 , 0 , n403 );
or_AQFP n404_( clk_6 , n402 , n403 , 0 , 0 , n404 );
and_AQFP n405_( clk_2 , splittern115ton370n405 , splittern396ton397n409 , 0 , 0 , n405 );
and_AQFP n406_( clk_4 , splitterG27ton406n407 , splitterfromn405 , 0 , 1 , n406 );
and_AQFP n407_( clk_4 , splitterG27ton406n407 , splitterfromn405 , 1 , 0 , n407 );
or_AQFP n408_( clk_6 , n406 , n407 , 0 , 0 , n408 );
and_AQFP n409_( clk_2 , splittern152ton374n409 , splittern396ton397n409 , 0 , 0 , n409 );
and_AQFP n410_( clk_4 , splitterG28ton410n411 , splitterfromn409 , 0 , 1 , n410 );
and_AQFP n411_( clk_4 , splitterG28ton410n411 , splitterfromn409 , 1 , 0 , n411 );
or_AQFP n412_( clk_6 , n410 , n411 , 0 , 0 , n412 );
and_AQFP n413_( clk_5 , splitterfromn250 , splittern272ton273n312 , 0 , 0 , n413 );
and_AQFP n414_( clk_6 , splittern359ton360n414 , n413 , 0 , 0 , n414 );
and_AQFP n415_( clk_8 , splittern172ton380n397 , splittern414ton415n427 , 0 , 0 , n415 );
or_AQFP n416_( clk_2 , splitterG29ton416n417 , splitterfromn415 , 0 , 0 , n416 );
and_AQFP n417_( clk_2 , splitterG29ton416n417 , splitterfromn415 , 0 , 0 , n417 );
and_AQFP n418_( clk_4 , n416 , n417 , 0 , 1 , n418 );
and_AQFP n419_( clk_8 , splittern191ton384n401 , splittern414ton415n427 , 0 , 0 , n419 );
and_AQFP n420_( clk_2 , splitterG30ton420n421 , splitterfromn419 , 0 , 1 , n420 );
and_AQFP n421_( clk_2 , splitterG30ton420n421 , splitterfromn419 , 1 , 0 , n421 );
or_AQFP n422_( clk_4 , n420 , n421 , 0 , 0 , n422 );
and_AQFP n423_( clk_8 , splittern115ton388n405 , splittern414ton415n427 , 0 , 0 , n423 );
and_AQFP n424_( clk_2 , splitterG31ton424n425 , splitterfromn423 , 0 , 1 , n424 );
and_AQFP n425_( clk_2 , splitterG31ton424n425 , splitterfromn423 , 1 , 0 , n425 );
or_AQFP n426_( clk_4 , n424 , n425 , 0 , 0 , n426 );
and_AQFP n427_( clk_8 , splittern152ton392n409 , splittern414ton415n427 , 0 , 0 , n427 );
or_AQFP n428_( clk_2 , splitterG32ton428n429 , splitterfromn427 , 0 , 0 , n428 );
and_AQFP n429_( clk_2 , splitterG32ton428n429 , splitterfromn427 , 0 , 0 , n429 );
and_AQFP n430_( clk_4 , n428 , n429 , 0 , 1 , n430 );
PO_AQFP G1324_( clk_8 , n285 , 1 , G1324 );
PO_AQFP G1325_( clk_8 , n289 , 1 , G1325 );
PO_AQFP G1326_( clk_8 , n293 , 1 , G1326 );
PO_AQFP G1327_( clk_8 , n297 , 1 , G1327 );
PO_AQFP G1328_( clk_8 , n303 , 1 , G1328 );
PO_AQFP G1329_( clk_8 , n307 , 1 , G1329 );
PO_AQFP G1330_( clk_8 , n311 , 1 , G1330 );
PO_AQFP G1331_( clk_8 , n315 , 1 , G1331 );
PO_AQFP G1332_( clk_8 , n322 , 1 , G1332 );
PO_AQFP G1333_( clk_8 , n326 , 1 , G1333 );
PO_AQFP G1334_( clk_8 , n330 , 1 , G1334 );
PO_AQFP G1335_( clk_8 , n334 , 1 , G1335 );
PO_AQFP G1336_( clk_8 , n340 , 1 , G1336 );
PO_AQFP G1337_( clk_8 , n344 , 1 , G1337 );
PO_AQFP G1338_( clk_8 , n348 , 1 , G1338 );
PO_AQFP G1339_( clk_8 , n352 , 1 , G1339 );
PO_AQFP G1340_( clk_8 , n365 , 1 , G1340 );
PO_AQFP G1341_( clk_8 , n369 , 1 , G1341 );
PO_AQFP G1342_( clk_8 , n373 , 1 , G1342 );
PO_AQFP G1343_( clk_8 , n377 , 1 , G1343 );
PO_AQFP G1344_( clk_8 , buf_n383_G1344_1 , 1 , G1344 );
PO_AQFP G1345_( clk_8 , buf_n387_G1345_1 , 1 , G1345 );
PO_AQFP G1346_( clk_8 , buf_n391_G1346_1 , 1 , G1346 );
PO_AQFP G1347_( clk_8 , buf_n395_G1347_1 , 1 , G1347 );
PO_AQFP G1348_( clk_8 , n400 , 1 , G1348 );
PO_AQFP G1349_( clk_8 , n404 , 1 , G1349 );
PO_AQFP G1350_( clk_8 , n408 , 1 , G1350 );
PO_AQFP G1351_( clk_8 , n412 , 1 , G1351 );
PO_AQFP G1352_( clk_8 , buf_n418_G1352_1 , 1 , G1352 );
PO_AQFP G1353_( clk_8 , buf_n422_G1353_1 , 1 , G1353 );
PO_AQFP G1354_( clk_8 , buf_n426_G1354_1 , 1 , G1354 );
PO_AQFP G1355_( clk_8 , buf_n430_G1355_1 , 1 , G1355 );
buf_AQFP buf_G33_n42_1_( clk_3 , G33 , 0 , buf_G33_n42_1 );
buf_AQFP buf_G34_n193_1_( clk_3 , G34 , 0 , buf_G34_n193_1 );
buf_AQFP buf_G35_n231_1_( clk_3 , G35 , 0 , buf_G35_n231_1 );
buf_AQFP buf_G36_n254_1_( clk_3 , G36 , 0 , buf_G36_n254_1 );
buf_AQFP buf_G37_n154_1_( clk_3 , G37 , 0 , buf_G37_n154_1 );
buf_AQFP buf_G39_n88_1_( clk_3 , G39 , 0 , buf_G39_n88_1 );
buf_AQFP buf_G40_n125_1_( clk_3 , G40 , 0 , buf_G40_n125_1 );
buf_AQFP buf_n42_splitterfromn42_1_( clk_7 , n42 , 0 , buf_n42_splitterfromn42_1 );
buf_AQFP buf_n88_splitterfromn88_1_( clk_7 , n88 , 0 , buf_n88_splitterfromn88_1 );
buf_AQFP buf_n125_splitterfromn125_1_( clk_6 , n125 , 0 , buf_n125_splitterfromn125_1 );
buf_AQFP buf_n154_splitterfromn154_1_( clk_6 , n154 , 0 , buf_n154_splitterfromn154_1 );
buf_AQFP buf_n173_splitterfromn173_2_( clk_5 , n173 , 0 , buf_n173_splitterfromn173_2 );
buf_AQFP buf_n173_splitterfromn173_1_( clk_7 , buf_n173_splitterfromn173_2 , 0 , buf_n173_splitterfromn173_1 );
buf_AQFP buf_n193_splitterfromn193_1_( clk_6 , n193 , 0 , buf_n193_splitterfromn193_1 );
buf_AQFP buf_n231_splitterfromn231_1_( clk_7 , n231 , 0 , buf_n231_splitterfromn231_1 );
buf_AQFP buf_n254_splitterfromn254_1_( clk_7 , n254 , 0 , buf_n254_splitterfromn254_1 );
buf_AQFP buf_n383_G1344_1_( clk_6 , n383 , 0 , buf_n383_G1344_1 );
buf_AQFP buf_n387_G1345_1_( clk_6 , n387 , 0 , buf_n387_G1345_1 );
buf_AQFP buf_n391_G1346_1_( clk_6 , n391 , 0 , buf_n391_G1346_1 );
buf_AQFP buf_n395_G1347_1_( clk_6 , n395 , 0 , buf_n395_G1347_1 );
buf_AQFP buf_n418_G1352_1_( clk_6 , n418 , 0 , buf_n418_G1352_1 );
buf_AQFP buf_n422_G1353_1_( clk_6 , n422 , 0 , buf_n422_G1353_1 );
buf_AQFP buf_n426_G1354_1_( clk_6 , n426 , 0 , buf_n426_G1354_1 );
buf_AQFP buf_n430_G1355_1_( clk_6 , n430 , 0 , buf_n430_G1355_1 );
buf_AQFP buf_splitterG1ton83n284_splitterG1ton283n284_12_( clk_5 , splitterG1ton83n284 , 0 , buf_splitterG1ton83n284_splitterG1ton283n284_12 );
buf_AQFP buf_splitterG1ton83n284_splitterG1ton283n284_11_( clk_7 , buf_splitterG1ton83n284_splitterG1ton283n284_12 , 0 , buf_splitterG1ton83n284_splitterG1ton283n284_11 );
buf_AQFP buf_splitterG1ton83n284_splitterG1ton283n284_10_( clk_1 , buf_splitterG1ton83n284_splitterG1ton283n284_11 , 0 , buf_splitterG1ton83n284_splitterG1ton283n284_10 );
buf_AQFP buf_splitterG1ton83n284_splitterG1ton283n284_9_( clk_3 , buf_splitterG1ton83n284_splitterG1ton283n284_10 , 0 , buf_splitterG1ton83n284_splitterG1ton283n284_9 );
buf_AQFP buf_splitterG1ton83n284_splitterG1ton283n284_8_( clk_5 , buf_splitterG1ton83n284_splitterG1ton283n284_9 , 0 , buf_splitterG1ton83n284_splitterG1ton283n284_8 );
buf_AQFP buf_splitterG1ton83n284_splitterG1ton283n284_7_( clk_7 , buf_splitterG1ton83n284_splitterG1ton283n284_8 , 0 , buf_splitterG1ton83n284_splitterG1ton283n284_7 );
buf_AQFP buf_splitterG1ton83n284_splitterG1ton283n284_6_( clk_1 , buf_splitterG1ton83n284_splitterG1ton283n284_7 , 0 , buf_splitterG1ton83n284_splitterG1ton283n284_6 );
buf_AQFP buf_splitterG1ton83n284_splitterG1ton283n284_5_( clk_3 , buf_splitterG1ton83n284_splitterG1ton283n284_6 , 0 , buf_splitterG1ton83n284_splitterG1ton283n284_5 );
buf_AQFP buf_splitterG1ton83n284_splitterG1ton283n284_4_( clk_5 , buf_splitterG1ton83n284_splitterG1ton283n284_5 , 0 , buf_splitterG1ton83n284_splitterG1ton283n284_4 );
buf_AQFP buf_splitterG1ton83n284_splitterG1ton283n284_3_( clk_7 , buf_splitterG1ton83n284_splitterG1ton283n284_4 , 0 , buf_splitterG1ton83n284_splitterG1ton283n284_3 );
buf_AQFP buf_splitterG1ton83n284_splitterG1ton283n284_2_( clk_1 , buf_splitterG1ton83n284_splitterG1ton283n284_3 , 0 , buf_splitterG1ton83n284_splitterG1ton283n284_2 );
buf_AQFP buf_splitterG1ton83n284_splitterG1ton283n284_1_( clk_3 , buf_splitterG1ton83n284_splitterG1ton283n284_2 , 0 , buf_splitterG1ton83n284_splitterG1ton283n284_1 );
buf_AQFP buf_splitterG10ton219n325_splitterG10ton324n325_11_( clk_5 , splitterG10ton219n325 , 0 , buf_splitterG10ton219n325_splitterG10ton324n325_11 );
buf_AQFP buf_splitterG10ton219n325_splitterG10ton324n325_10_( clk_7 , buf_splitterG10ton219n325_splitterG10ton324n325_11 , 0 , buf_splitterG10ton219n325_splitterG10ton324n325_10 );
buf_AQFP buf_splitterG10ton219n325_splitterG10ton324n325_9_( clk_1 , buf_splitterG10ton219n325_splitterG10ton324n325_10 , 0 , buf_splitterG10ton219n325_splitterG10ton324n325_9 );
buf_AQFP buf_splitterG10ton219n325_splitterG10ton324n325_8_( clk_3 , buf_splitterG10ton219n325_splitterG10ton324n325_9 , 0 , buf_splitterG10ton219n325_splitterG10ton324n325_8 );
buf_AQFP buf_splitterG10ton219n325_splitterG10ton324n325_7_( clk_5 , buf_splitterG10ton219n325_splitterG10ton324n325_8 , 0 , buf_splitterG10ton219n325_splitterG10ton324n325_7 );
buf_AQFP buf_splitterG10ton219n325_splitterG10ton324n325_6_( clk_7 , buf_splitterG10ton219n325_splitterG10ton324n325_7 , 0 , buf_splitterG10ton219n325_splitterG10ton324n325_6 );
buf_AQFP buf_splitterG10ton219n325_splitterG10ton324n325_5_( clk_1 , buf_splitterG10ton219n325_splitterG10ton324n325_6 , 0 , buf_splitterG10ton219n325_splitterG10ton324n325_5 );
buf_AQFP buf_splitterG10ton219n325_splitterG10ton324n325_4_( clk_3 , buf_splitterG10ton219n325_splitterG10ton324n325_5 , 0 , buf_splitterG10ton219n325_splitterG10ton324n325_4 );
buf_AQFP buf_splitterG10ton219n325_splitterG10ton324n325_3_( clk_5 , buf_splitterG10ton219n325_splitterG10ton324n325_4 , 0 , buf_splitterG10ton219n325_splitterG10ton324n325_3 );
buf_AQFP buf_splitterG10ton219n325_splitterG10ton324n325_2_( clk_7 , buf_splitterG10ton219n325_splitterG10ton324n325_3 , 0 , buf_splitterG10ton219n325_splitterG10ton324n325_2 );
buf_AQFP buf_splitterG10ton219n325_splitterG10ton324n325_1_( clk_1 , buf_splitterG10ton219n325_splitterG10ton324n325_2 , 0 , buf_splitterG10ton219n325_splitterG10ton324n325_1 );
buf_AQFP buf_splitterG11ton235n329_splitterG11ton328n329_11_( clk_5 , splitterG11ton235n329 , 0 , buf_splitterG11ton235n329_splitterG11ton328n329_11 );
buf_AQFP buf_splitterG11ton235n329_splitterG11ton328n329_10_( clk_7 , buf_splitterG11ton235n329_splitterG11ton328n329_11 , 0 , buf_splitterG11ton235n329_splitterG11ton328n329_10 );
buf_AQFP buf_splitterG11ton235n329_splitterG11ton328n329_9_( clk_1 , buf_splitterG11ton235n329_splitterG11ton328n329_10 , 0 , buf_splitterG11ton235n329_splitterG11ton328n329_9 );
buf_AQFP buf_splitterG11ton235n329_splitterG11ton328n329_8_( clk_3 , buf_splitterG11ton235n329_splitterG11ton328n329_9 , 0 , buf_splitterG11ton235n329_splitterG11ton328n329_8 );
buf_AQFP buf_splitterG11ton235n329_splitterG11ton328n329_7_( clk_5 , buf_splitterG11ton235n329_splitterG11ton328n329_8 , 0 , buf_splitterG11ton235n329_splitterG11ton328n329_7 );
buf_AQFP buf_splitterG11ton235n329_splitterG11ton328n329_6_( clk_7 , buf_splitterG11ton235n329_splitterG11ton328n329_7 , 0 , buf_splitterG11ton235n329_splitterG11ton328n329_6 );
buf_AQFP buf_splitterG11ton235n329_splitterG11ton328n329_5_( clk_1 , buf_splitterG11ton235n329_splitterG11ton328n329_6 , 0 , buf_splitterG11ton235n329_splitterG11ton328n329_5 );
buf_AQFP buf_splitterG11ton235n329_splitterG11ton328n329_4_( clk_3 , buf_splitterG11ton235n329_splitterG11ton328n329_5 , 0 , buf_splitterG11ton235n329_splitterG11ton328n329_4 );
buf_AQFP buf_splitterG11ton235n329_splitterG11ton328n329_3_( clk_5 , buf_splitterG11ton235n329_splitterG11ton328n329_4 , 0 , buf_splitterG11ton235n329_splitterG11ton328n329_3 );
buf_AQFP buf_splitterG11ton235n329_splitterG11ton328n329_2_( clk_7 , buf_splitterG11ton235n329_splitterG11ton328n329_3 , 0 , buf_splitterG11ton235n329_splitterG11ton328n329_2 );
buf_AQFP buf_splitterG11ton235n329_splitterG11ton328n329_1_( clk_1 , buf_splitterG11ton235n329_splitterG11ton328n329_2 , 0 , buf_splitterG11ton235n329_splitterG11ton328n329_1 );
buf_AQFP buf_splitterG12ton93n333_splitterG12ton332n333_11_( clk_5 , splitterG12ton93n333 , 0 , buf_splitterG12ton93n333_splitterG12ton332n333_11 );
buf_AQFP buf_splitterG12ton93n333_splitterG12ton332n333_10_( clk_7 , buf_splitterG12ton93n333_splitterG12ton332n333_11 , 0 , buf_splitterG12ton93n333_splitterG12ton332n333_10 );
buf_AQFP buf_splitterG12ton93n333_splitterG12ton332n333_9_( clk_1 , buf_splitterG12ton93n333_splitterG12ton332n333_10 , 0 , buf_splitterG12ton93n333_splitterG12ton332n333_9 );
buf_AQFP buf_splitterG12ton93n333_splitterG12ton332n333_8_( clk_3 , buf_splitterG12ton93n333_splitterG12ton332n333_9 , 0 , buf_splitterG12ton93n333_splitterG12ton332n333_8 );
buf_AQFP buf_splitterG12ton93n333_splitterG12ton332n333_7_( clk_5 , buf_splitterG12ton93n333_splitterG12ton332n333_8 , 0 , buf_splitterG12ton93n333_splitterG12ton332n333_7 );
buf_AQFP buf_splitterG12ton93n333_splitterG12ton332n333_6_( clk_7 , buf_splitterG12ton93n333_splitterG12ton332n333_7 , 0 , buf_splitterG12ton93n333_splitterG12ton332n333_6 );
buf_AQFP buf_splitterG12ton93n333_splitterG12ton332n333_5_( clk_1 , buf_splitterG12ton93n333_splitterG12ton332n333_6 , 0 , buf_splitterG12ton93n333_splitterG12ton332n333_5 );
buf_AQFP buf_splitterG12ton93n333_splitterG12ton332n333_4_( clk_3 , buf_splitterG12ton93n333_splitterG12ton332n333_5 , 0 , buf_splitterG12ton93n333_splitterG12ton332n333_4 );
buf_AQFP buf_splitterG12ton93n333_splitterG12ton332n333_3_( clk_5 , buf_splitterG12ton93n333_splitterG12ton332n333_4 , 0 , buf_splitterG12ton93n333_splitterG12ton332n333_3 );
buf_AQFP buf_splitterG12ton93n333_splitterG12ton332n333_2_( clk_7 , buf_splitterG12ton93n333_splitterG12ton332n333_3 , 0 , buf_splitterG12ton93n333_splitterG12ton332n333_2 );
buf_AQFP buf_splitterG12ton93n333_splitterG12ton332n333_1_( clk_1 , buf_splitterG12ton93n333_splitterG12ton332n333_2 , 0 , buf_splitterG12ton93n333_splitterG12ton332n333_1 );
buf_AQFP buf_splitterG13ton65n339_splitterG13ton338n339_11_( clk_5 , splitterG13ton65n339 , 0 , buf_splitterG13ton65n339_splitterG13ton338n339_11 );
buf_AQFP buf_splitterG13ton65n339_splitterG13ton338n339_10_( clk_7 , buf_splitterG13ton65n339_splitterG13ton338n339_11 , 0 , buf_splitterG13ton65n339_splitterG13ton338n339_10 );
buf_AQFP buf_splitterG13ton65n339_splitterG13ton338n339_9_( clk_1 , buf_splitterG13ton65n339_splitterG13ton338n339_10 , 0 , buf_splitterG13ton65n339_splitterG13ton338n339_9 );
buf_AQFP buf_splitterG13ton65n339_splitterG13ton338n339_8_( clk_3 , buf_splitterG13ton65n339_splitterG13ton338n339_9 , 0 , buf_splitterG13ton65n339_splitterG13ton338n339_8 );
buf_AQFP buf_splitterG13ton65n339_splitterG13ton338n339_7_( clk_5 , buf_splitterG13ton65n339_splitterG13ton338n339_8 , 0 , buf_splitterG13ton65n339_splitterG13ton338n339_7 );
buf_AQFP buf_splitterG13ton65n339_splitterG13ton338n339_6_( clk_7 , buf_splitterG13ton65n339_splitterG13ton338n339_7 , 0 , buf_splitterG13ton65n339_splitterG13ton338n339_6 );
buf_AQFP buf_splitterG13ton65n339_splitterG13ton338n339_5_( clk_1 , buf_splitterG13ton65n339_splitterG13ton338n339_6 , 0 , buf_splitterG13ton65n339_splitterG13ton338n339_5 );
buf_AQFP buf_splitterG13ton65n339_splitterG13ton338n339_4_( clk_3 , buf_splitterG13ton65n339_splitterG13ton338n339_5 , 0 , buf_splitterG13ton65n339_splitterG13ton338n339_4 );
buf_AQFP buf_splitterG13ton65n339_splitterG13ton338n339_3_( clk_5 , buf_splitterG13ton65n339_splitterG13ton338n339_4 , 0 , buf_splitterG13ton65n339_splitterG13ton338n339_3 );
buf_AQFP buf_splitterG13ton65n339_splitterG13ton338n339_2_( clk_7 , buf_splitterG13ton65n339_splitterG13ton338n339_3 , 0 , buf_splitterG13ton65n339_splitterG13ton338n339_2 );
buf_AQFP buf_splitterG13ton65n339_splitterG13ton338n339_1_( clk_1 , buf_splitterG13ton65n339_splitterG13ton338n339_2 , 0 , buf_splitterG13ton65n339_splitterG13ton338n339_1 );
buf_AQFP buf_splitterG14ton216n343_splitterG14ton342n343_11_( clk_5 , splitterG14ton216n343 , 0 , buf_splitterG14ton216n343_splitterG14ton342n343_11 );
buf_AQFP buf_splitterG14ton216n343_splitterG14ton342n343_10_( clk_7 , buf_splitterG14ton216n343_splitterG14ton342n343_11 , 0 , buf_splitterG14ton216n343_splitterG14ton342n343_10 );
buf_AQFP buf_splitterG14ton216n343_splitterG14ton342n343_9_( clk_1 , buf_splitterG14ton216n343_splitterG14ton342n343_10 , 0 , buf_splitterG14ton216n343_splitterG14ton342n343_9 );
buf_AQFP buf_splitterG14ton216n343_splitterG14ton342n343_8_( clk_3 , buf_splitterG14ton216n343_splitterG14ton342n343_9 , 0 , buf_splitterG14ton216n343_splitterG14ton342n343_8 );
buf_AQFP buf_splitterG14ton216n343_splitterG14ton342n343_7_( clk_5 , buf_splitterG14ton216n343_splitterG14ton342n343_8 , 0 , buf_splitterG14ton216n343_splitterG14ton342n343_7 );
buf_AQFP buf_splitterG14ton216n343_splitterG14ton342n343_6_( clk_7 , buf_splitterG14ton216n343_splitterG14ton342n343_7 , 0 , buf_splitterG14ton216n343_splitterG14ton342n343_6 );
buf_AQFP buf_splitterG14ton216n343_splitterG14ton342n343_5_( clk_1 , buf_splitterG14ton216n343_splitterG14ton342n343_6 , 0 , buf_splitterG14ton216n343_splitterG14ton342n343_5 );
buf_AQFP buf_splitterG14ton216n343_splitterG14ton342n343_4_( clk_3 , buf_splitterG14ton216n343_splitterG14ton342n343_5 , 0 , buf_splitterG14ton216n343_splitterG14ton342n343_4 );
buf_AQFP buf_splitterG14ton216n343_splitterG14ton342n343_3_( clk_5 , buf_splitterG14ton216n343_splitterG14ton342n343_4 , 0 , buf_splitterG14ton216n343_splitterG14ton342n343_3 );
buf_AQFP buf_splitterG14ton216n343_splitterG14ton342n343_2_( clk_7 , buf_splitterG14ton216n343_splitterG14ton342n343_3 , 0 , buf_splitterG14ton216n343_splitterG14ton342n343_2 );
buf_AQFP buf_splitterG14ton216n343_splitterG14ton342n343_1_( clk_1 , buf_splitterG14ton216n343_splitterG14ton342n343_2 , 0 , buf_splitterG14ton216n343_splitterG14ton342n343_1 );
buf_AQFP buf_splitterG15ton236n347_splitterG15ton346n347_10_( clk_6 , splitterG15ton236n347 , 0 , buf_splitterG15ton236n347_splitterG15ton346n347_10 );
buf_AQFP buf_splitterG15ton236n347_splitterG15ton346n347_9_( clk_8 , buf_splitterG15ton236n347_splitterG15ton346n347_10 , 0 , buf_splitterG15ton236n347_splitterG15ton346n347_9 );
buf_AQFP buf_splitterG15ton236n347_splitterG15ton346n347_8_( clk_2 , buf_splitterG15ton236n347_splitterG15ton346n347_9 , 0 , buf_splitterG15ton236n347_splitterG15ton346n347_8 );
buf_AQFP buf_splitterG15ton236n347_splitterG15ton346n347_7_( clk_4 , buf_splitterG15ton236n347_splitterG15ton346n347_8 , 0 , buf_splitterG15ton236n347_splitterG15ton346n347_7 );
buf_AQFP buf_splitterG15ton236n347_splitterG15ton346n347_6_( clk_6 , buf_splitterG15ton236n347_splitterG15ton346n347_7 , 0 , buf_splitterG15ton236n347_splitterG15ton346n347_6 );
buf_AQFP buf_splitterG15ton236n347_splitterG15ton346n347_5_( clk_8 , buf_splitterG15ton236n347_splitterG15ton346n347_6 , 0 , buf_splitterG15ton236n347_splitterG15ton346n347_5 );
buf_AQFP buf_splitterG15ton236n347_splitterG15ton346n347_4_( clk_2 , buf_splitterG15ton236n347_splitterG15ton346n347_5 , 0 , buf_splitterG15ton236n347_splitterG15ton346n347_4 );
buf_AQFP buf_splitterG15ton236n347_splitterG15ton346n347_3_( clk_4 , buf_splitterG15ton236n347_splitterG15ton346n347_4 , 0 , buf_splitterG15ton236n347_splitterG15ton346n347_3 );
buf_AQFP buf_splitterG15ton236n347_splitterG15ton346n347_2_( clk_6 , buf_splitterG15ton236n347_splitterG15ton346n347_3 , 0 , buf_splitterG15ton236n347_splitterG15ton346n347_2 );
buf_AQFP buf_splitterG15ton236n347_splitterG15ton346n347_1_( clk_8 , buf_splitterG15ton236n347_splitterG15ton346n347_2 , 0 , buf_splitterG15ton236n347_splitterG15ton346n347_1 );
buf_AQFP buf_splitterG16ton262n351_splitterG16ton350n351_10_( clk_6 , splitterG16ton262n351 , 0 , buf_splitterG16ton262n351_splitterG16ton350n351_10 );
buf_AQFP buf_splitterG16ton262n351_splitterG16ton350n351_9_( clk_8 , buf_splitterG16ton262n351_splitterG16ton350n351_10 , 0 , buf_splitterG16ton262n351_splitterG16ton350n351_9 );
buf_AQFP buf_splitterG16ton262n351_splitterG16ton350n351_8_( clk_2 , buf_splitterG16ton262n351_splitterG16ton350n351_9 , 0 , buf_splitterG16ton262n351_splitterG16ton350n351_8 );
buf_AQFP buf_splitterG16ton262n351_splitterG16ton350n351_7_( clk_4 , buf_splitterG16ton262n351_splitterG16ton350n351_8 , 0 , buf_splitterG16ton262n351_splitterG16ton350n351_7 );
buf_AQFP buf_splitterG16ton262n351_splitterG16ton350n351_6_( clk_6 , buf_splitterG16ton262n351_splitterG16ton350n351_7 , 0 , buf_splitterG16ton262n351_splitterG16ton350n351_6 );
buf_AQFP buf_splitterG16ton262n351_splitterG16ton350n351_5_( clk_8 , buf_splitterG16ton262n351_splitterG16ton350n351_6 , 0 , buf_splitterG16ton262n351_splitterG16ton350n351_5 );
buf_AQFP buf_splitterG16ton262n351_splitterG16ton350n351_4_( clk_2 , buf_splitterG16ton262n351_splitterG16ton350n351_5 , 0 , buf_splitterG16ton262n351_splitterG16ton350n351_4 );
buf_AQFP buf_splitterG16ton262n351_splitterG16ton350n351_3_( clk_4 , buf_splitterG16ton262n351_splitterG16ton350n351_4 , 0 , buf_splitterG16ton262n351_splitterG16ton350n351_3 );
buf_AQFP buf_splitterG16ton262n351_splitterG16ton350n351_2_( clk_6 , buf_splitterG16ton262n351_splitterG16ton350n351_3 , 0 , buf_splitterG16ton262n351_splitterG16ton350n351_2 );
buf_AQFP buf_splitterG16ton262n351_splitterG16ton350n351_1_( clk_8 , buf_splitterG16ton262n351_splitterG16ton350n351_2 , 0 , buf_splitterG16ton262n351_splitterG16ton350n351_1 );
buf_AQFP buf_splitterG17ton44n364_splitterG17ton363n364_11_( clk_5 , splitterG17ton44n364 , 0 , buf_splitterG17ton44n364_splitterG17ton363n364_11 );
buf_AQFP buf_splitterG17ton44n364_splitterG17ton363n364_10_( clk_7 , buf_splitterG17ton44n364_splitterG17ton363n364_11 , 0 , buf_splitterG17ton44n364_splitterG17ton363n364_10 );
buf_AQFP buf_splitterG17ton44n364_splitterG17ton363n364_9_( clk_1 , buf_splitterG17ton44n364_splitterG17ton363n364_10 , 0 , buf_splitterG17ton44n364_splitterG17ton363n364_9 );
buf_AQFP buf_splitterG17ton44n364_splitterG17ton363n364_8_( clk_3 , buf_splitterG17ton44n364_splitterG17ton363n364_9 , 0 , buf_splitterG17ton44n364_splitterG17ton363n364_8 );
buf_AQFP buf_splitterG17ton44n364_splitterG17ton363n364_7_( clk_5 , buf_splitterG17ton44n364_splitterG17ton363n364_8 , 0 , buf_splitterG17ton44n364_splitterG17ton363n364_7 );
buf_AQFP buf_splitterG17ton44n364_splitterG17ton363n364_6_( clk_7 , buf_splitterG17ton44n364_splitterG17ton363n364_7 , 0 , buf_splitterG17ton44n364_splitterG17ton363n364_6 );
buf_AQFP buf_splitterG17ton44n364_splitterG17ton363n364_5_( clk_1 , buf_splitterG17ton44n364_splitterG17ton363n364_6 , 0 , buf_splitterG17ton44n364_splitterG17ton363n364_5 );
buf_AQFP buf_splitterG17ton44n364_splitterG17ton363n364_4_( clk_3 , buf_splitterG17ton44n364_splitterG17ton363n364_5 , 0 , buf_splitterG17ton44n364_splitterG17ton363n364_4 );
buf_AQFP buf_splitterG17ton44n364_splitterG17ton363n364_3_( clk_5 , buf_splitterG17ton44n364_splitterG17ton363n364_4 , 0 , buf_splitterG17ton44n364_splitterG17ton363n364_3 );
buf_AQFP buf_splitterG17ton44n364_splitterG17ton363n364_2_( clk_7 , buf_splitterG17ton44n364_splitterG17ton363n364_3 , 0 , buf_splitterG17ton44n364_splitterG17ton363n364_2 );
buf_AQFP buf_splitterG17ton44n364_splitterG17ton363n364_1_( clk_1 , buf_splitterG17ton44n364_splitterG17ton363n364_2 , 0 , buf_splitterG17ton44n364_splitterG17ton363n364_1 );
buf_AQFP buf_splitterG18ton47n368_splitterG18ton367n368_11_( clk_5 , splitterG18ton47n368 , 0 , buf_splitterG18ton47n368_splitterG18ton367n368_11 );
buf_AQFP buf_splitterG18ton47n368_splitterG18ton367n368_10_( clk_7 , buf_splitterG18ton47n368_splitterG18ton367n368_11 , 0 , buf_splitterG18ton47n368_splitterG18ton367n368_10 );
buf_AQFP buf_splitterG18ton47n368_splitterG18ton367n368_9_( clk_1 , buf_splitterG18ton47n368_splitterG18ton367n368_10 , 0 , buf_splitterG18ton47n368_splitterG18ton367n368_9 );
buf_AQFP buf_splitterG18ton47n368_splitterG18ton367n368_8_( clk_3 , buf_splitterG18ton47n368_splitterG18ton367n368_9 , 0 , buf_splitterG18ton47n368_splitterG18ton367n368_8 );
buf_AQFP buf_splitterG18ton47n368_splitterG18ton367n368_7_( clk_5 , buf_splitterG18ton47n368_splitterG18ton367n368_8 , 0 , buf_splitterG18ton47n368_splitterG18ton367n368_7 );
buf_AQFP buf_splitterG18ton47n368_splitterG18ton367n368_6_( clk_7 , buf_splitterG18ton47n368_splitterG18ton367n368_7 , 0 , buf_splitterG18ton47n368_splitterG18ton367n368_6 );
buf_AQFP buf_splitterG18ton47n368_splitterG18ton367n368_5_( clk_1 , buf_splitterG18ton47n368_splitterG18ton367n368_6 , 0 , buf_splitterG18ton47n368_splitterG18ton367n368_5 );
buf_AQFP buf_splitterG18ton47n368_splitterG18ton367n368_4_( clk_3 , buf_splitterG18ton47n368_splitterG18ton367n368_5 , 0 , buf_splitterG18ton47n368_splitterG18ton367n368_4 );
buf_AQFP buf_splitterG18ton47n368_splitterG18ton367n368_3_( clk_5 , buf_splitterG18ton47n368_splitterG18ton367n368_4 , 0 , buf_splitterG18ton47n368_splitterG18ton367n368_3 );
buf_AQFP buf_splitterG18ton47n368_splitterG18ton367n368_2_( clk_7 , buf_splitterG18ton47n368_splitterG18ton367n368_3 , 0 , buf_splitterG18ton47n368_splitterG18ton367n368_2 );
buf_AQFP buf_splitterG18ton47n368_splitterG18ton367n368_1_( clk_1 , buf_splitterG18ton47n368_splitterG18ton367n368_2 , 0 , buf_splitterG18ton47n368_splitterG18ton367n368_1 );
buf_AQFP buf_splitterG19ton44n372_splitterG19ton371n372_11_( clk_5 , splitterG19ton44n372 , 0 , buf_splitterG19ton44n372_splitterG19ton371n372_11 );
buf_AQFP buf_splitterG19ton44n372_splitterG19ton371n372_10_( clk_7 , buf_splitterG19ton44n372_splitterG19ton371n372_11 , 0 , buf_splitterG19ton44n372_splitterG19ton371n372_10 );
buf_AQFP buf_splitterG19ton44n372_splitterG19ton371n372_9_( clk_1 , buf_splitterG19ton44n372_splitterG19ton371n372_10 , 0 , buf_splitterG19ton44n372_splitterG19ton371n372_9 );
buf_AQFP buf_splitterG19ton44n372_splitterG19ton371n372_8_( clk_3 , buf_splitterG19ton44n372_splitterG19ton371n372_9 , 0 , buf_splitterG19ton44n372_splitterG19ton371n372_8 );
buf_AQFP buf_splitterG19ton44n372_splitterG19ton371n372_7_( clk_5 , buf_splitterG19ton44n372_splitterG19ton371n372_8 , 0 , buf_splitterG19ton44n372_splitterG19ton371n372_7 );
buf_AQFP buf_splitterG19ton44n372_splitterG19ton371n372_6_( clk_7 , buf_splitterG19ton44n372_splitterG19ton371n372_7 , 0 , buf_splitterG19ton44n372_splitterG19ton371n372_6 );
buf_AQFP buf_splitterG19ton44n372_splitterG19ton371n372_5_( clk_1 , buf_splitterG19ton44n372_splitterG19ton371n372_6 , 0 , buf_splitterG19ton44n372_splitterG19ton371n372_5 );
buf_AQFP buf_splitterG19ton44n372_splitterG19ton371n372_4_( clk_3 , buf_splitterG19ton44n372_splitterG19ton371n372_5 , 0 , buf_splitterG19ton44n372_splitterG19ton371n372_4 );
buf_AQFP buf_splitterG19ton44n372_splitterG19ton371n372_3_( clk_5 , buf_splitterG19ton44n372_splitterG19ton371n372_4 , 0 , buf_splitterG19ton44n372_splitterG19ton371n372_3 );
buf_AQFP buf_splitterG19ton44n372_splitterG19ton371n372_2_( clk_7 , buf_splitterG19ton44n372_splitterG19ton371n372_3 , 0 , buf_splitterG19ton44n372_splitterG19ton371n372_2 );
buf_AQFP buf_splitterG19ton44n372_splitterG19ton371n372_1_( clk_1 , buf_splitterG19ton44n372_splitterG19ton371n372_2 , 0 , buf_splitterG19ton44n372_splitterG19ton371n372_1 );
buf_AQFP buf_splitterG2ton216n288_splitterG2ton287n288_12_( clk_5 , splitterG2ton216n288 , 0 , buf_splitterG2ton216n288_splitterG2ton287n288_12 );
buf_AQFP buf_splitterG2ton216n288_splitterG2ton287n288_11_( clk_7 , buf_splitterG2ton216n288_splitterG2ton287n288_12 , 0 , buf_splitterG2ton216n288_splitterG2ton287n288_11 );
buf_AQFP buf_splitterG2ton216n288_splitterG2ton287n288_10_( clk_1 , buf_splitterG2ton216n288_splitterG2ton287n288_11 , 0 , buf_splitterG2ton216n288_splitterG2ton287n288_10 );
buf_AQFP buf_splitterG2ton216n288_splitterG2ton287n288_9_( clk_3 , buf_splitterG2ton216n288_splitterG2ton287n288_10 , 0 , buf_splitterG2ton216n288_splitterG2ton287n288_9 );
buf_AQFP buf_splitterG2ton216n288_splitterG2ton287n288_8_( clk_5 , buf_splitterG2ton216n288_splitterG2ton287n288_9 , 0 , buf_splitterG2ton216n288_splitterG2ton287n288_8 );
buf_AQFP buf_splitterG2ton216n288_splitterG2ton287n288_7_( clk_7 , buf_splitterG2ton216n288_splitterG2ton287n288_8 , 0 , buf_splitterG2ton216n288_splitterG2ton287n288_7 );
buf_AQFP buf_splitterG2ton216n288_splitterG2ton287n288_6_( clk_1 , buf_splitterG2ton216n288_splitterG2ton287n288_7 , 0 , buf_splitterG2ton216n288_splitterG2ton287n288_6 );
buf_AQFP buf_splitterG2ton216n288_splitterG2ton287n288_5_( clk_3 , buf_splitterG2ton216n288_splitterG2ton287n288_6 , 0 , buf_splitterG2ton216n288_splitterG2ton287n288_5 );
buf_AQFP buf_splitterG2ton216n288_splitterG2ton287n288_4_( clk_5 , buf_splitterG2ton216n288_splitterG2ton287n288_5 , 0 , buf_splitterG2ton216n288_splitterG2ton287n288_4 );
buf_AQFP buf_splitterG2ton216n288_splitterG2ton287n288_3_( clk_7 , buf_splitterG2ton216n288_splitterG2ton287n288_4 , 0 , buf_splitterG2ton216n288_splitterG2ton287n288_3 );
buf_AQFP buf_splitterG2ton216n288_splitterG2ton287n288_2_( clk_1 , buf_splitterG2ton216n288_splitterG2ton287n288_3 , 0 , buf_splitterG2ton216n288_splitterG2ton287n288_2 );
buf_AQFP buf_splitterG2ton216n288_splitterG2ton287n288_1_( clk_3 , buf_splitterG2ton216n288_splitterG2ton287n288_2 , 0 , buf_splitterG2ton216n288_splitterG2ton287n288_1 );
buf_AQFP buf_splitterG20ton47n376_splitterG20ton375n376_11_( clk_5 , splitterG20ton47n376 , 0 , buf_splitterG20ton47n376_splitterG20ton375n376_11 );
buf_AQFP buf_splitterG20ton47n376_splitterG20ton375n376_10_( clk_7 , buf_splitterG20ton47n376_splitterG20ton375n376_11 , 0 , buf_splitterG20ton47n376_splitterG20ton375n376_10 );
buf_AQFP buf_splitterG20ton47n376_splitterG20ton375n376_9_( clk_1 , buf_splitterG20ton47n376_splitterG20ton375n376_10 , 0 , buf_splitterG20ton47n376_splitterG20ton375n376_9 );
buf_AQFP buf_splitterG20ton47n376_splitterG20ton375n376_8_( clk_3 , buf_splitterG20ton47n376_splitterG20ton375n376_9 , 0 , buf_splitterG20ton47n376_splitterG20ton375n376_8 );
buf_AQFP buf_splitterG20ton47n376_splitterG20ton375n376_7_( clk_5 , buf_splitterG20ton47n376_splitterG20ton375n376_8 , 0 , buf_splitterG20ton47n376_splitterG20ton375n376_7 );
buf_AQFP buf_splitterG20ton47n376_splitterG20ton375n376_6_( clk_7 , buf_splitterG20ton47n376_splitterG20ton375n376_7 , 0 , buf_splitterG20ton47n376_splitterG20ton375n376_6 );
buf_AQFP buf_splitterG20ton47n376_splitterG20ton375n376_5_( clk_1 , buf_splitterG20ton47n376_splitterG20ton375n376_6 , 0 , buf_splitterG20ton47n376_splitterG20ton375n376_5 );
buf_AQFP buf_splitterG20ton47n376_splitterG20ton375n376_4_( clk_3 , buf_splitterG20ton47n376_splitterG20ton375n376_5 , 0 , buf_splitterG20ton47n376_splitterG20ton375n376_4 );
buf_AQFP buf_splitterG20ton47n376_splitterG20ton375n376_3_( clk_5 , buf_splitterG20ton47n376_splitterG20ton375n376_4 , 0 , buf_splitterG20ton47n376_splitterG20ton375n376_3 );
buf_AQFP buf_splitterG20ton47n376_splitterG20ton375n376_2_( clk_7 , buf_splitterG20ton47n376_splitterG20ton375n376_3 , 0 , buf_splitterG20ton47n376_splitterG20ton375n376_2 );
buf_AQFP buf_splitterG20ton47n376_splitterG20ton375n376_1_( clk_1 , buf_splitterG20ton47n376_splitterG20ton375n376_2 , 0 , buf_splitterG20ton47n376_splitterG20ton375n376_1 );
buf_AQFP buf_splitterG21ton59n382_splitterG21ton381n382_10_( clk_5 , splitterG21ton59n382 , 0 , buf_splitterG21ton59n382_splitterG21ton381n382_10 );
buf_AQFP buf_splitterG21ton59n382_splitterG21ton381n382_9_( clk_7 , buf_splitterG21ton59n382_splitterG21ton381n382_10 , 0 , buf_splitterG21ton59n382_splitterG21ton381n382_9 );
buf_AQFP buf_splitterG21ton59n382_splitterG21ton381n382_8_( clk_1 , buf_splitterG21ton59n382_splitterG21ton381n382_9 , 0 , buf_splitterG21ton59n382_splitterG21ton381n382_8 );
buf_AQFP buf_splitterG21ton59n382_splitterG21ton381n382_7_( clk_3 , buf_splitterG21ton59n382_splitterG21ton381n382_8 , 0 , buf_splitterG21ton59n382_splitterG21ton381n382_7 );
buf_AQFP buf_splitterG21ton59n382_splitterG21ton381n382_6_( clk_5 , buf_splitterG21ton59n382_splitterG21ton381n382_7 , 0 , buf_splitterG21ton59n382_splitterG21ton381n382_6 );
buf_AQFP buf_splitterG21ton59n382_splitterG21ton381n382_5_( clk_7 , buf_splitterG21ton59n382_splitterG21ton381n382_6 , 0 , buf_splitterG21ton59n382_splitterG21ton381n382_5 );
buf_AQFP buf_splitterG21ton59n382_splitterG21ton381n382_4_( clk_1 , buf_splitterG21ton59n382_splitterG21ton381n382_5 , 0 , buf_splitterG21ton59n382_splitterG21ton381n382_4 );
buf_AQFP buf_splitterG21ton59n382_splitterG21ton381n382_3_( clk_3 , buf_splitterG21ton59n382_splitterG21ton381n382_4 , 0 , buf_splitterG21ton59n382_splitterG21ton381n382_3 );
buf_AQFP buf_splitterG21ton59n382_splitterG21ton381n382_2_( clk_5 , buf_splitterG21ton59n382_splitterG21ton381n382_3 , 0 , buf_splitterG21ton59n382_splitterG21ton381n382_2 );
buf_AQFP buf_splitterG21ton59n382_splitterG21ton381n382_1_( clk_7 , buf_splitterG21ton59n382_splitterG21ton381n382_2 , 0 , buf_splitterG21ton59n382_splitterG21ton381n382_1 );
buf_AQFP buf_splitterG22ton56n386_splitterG22ton385n386_10_( clk_5 , splitterG22ton56n386 , 0 , buf_splitterG22ton56n386_splitterG22ton385n386_10 );
buf_AQFP buf_splitterG22ton56n386_splitterG22ton385n386_9_( clk_7 , buf_splitterG22ton56n386_splitterG22ton385n386_10 , 0 , buf_splitterG22ton56n386_splitterG22ton385n386_9 );
buf_AQFP buf_splitterG22ton56n386_splitterG22ton385n386_8_( clk_1 , buf_splitterG22ton56n386_splitterG22ton385n386_9 , 0 , buf_splitterG22ton56n386_splitterG22ton385n386_8 );
buf_AQFP buf_splitterG22ton56n386_splitterG22ton385n386_7_( clk_3 , buf_splitterG22ton56n386_splitterG22ton385n386_8 , 0 , buf_splitterG22ton56n386_splitterG22ton385n386_7 );
buf_AQFP buf_splitterG22ton56n386_splitterG22ton385n386_6_( clk_5 , buf_splitterG22ton56n386_splitterG22ton385n386_7 , 0 , buf_splitterG22ton56n386_splitterG22ton385n386_6 );
buf_AQFP buf_splitterG22ton56n386_splitterG22ton385n386_5_( clk_7 , buf_splitterG22ton56n386_splitterG22ton385n386_6 , 0 , buf_splitterG22ton56n386_splitterG22ton385n386_5 );
buf_AQFP buf_splitterG22ton56n386_splitterG22ton385n386_4_( clk_1 , buf_splitterG22ton56n386_splitterG22ton385n386_5 , 0 , buf_splitterG22ton56n386_splitterG22ton385n386_4 );
buf_AQFP buf_splitterG22ton56n386_splitterG22ton385n386_3_( clk_3 , buf_splitterG22ton56n386_splitterG22ton385n386_4 , 0 , buf_splitterG22ton56n386_splitterG22ton385n386_3 );
buf_AQFP buf_splitterG22ton56n386_splitterG22ton385n386_2_( clk_5 , buf_splitterG22ton56n386_splitterG22ton385n386_3 , 0 , buf_splitterG22ton56n386_splitterG22ton385n386_2 );
buf_AQFP buf_splitterG22ton56n386_splitterG22ton385n386_1_( clk_7 , buf_splitterG22ton56n386_splitterG22ton385n386_2 , 0 , buf_splitterG22ton56n386_splitterG22ton385n386_1 );
buf_AQFP buf_splitterG23ton56n390_splitterG23ton389n390_10_( clk_5 , splitterG23ton56n390 , 0 , buf_splitterG23ton56n390_splitterG23ton389n390_10 );
buf_AQFP buf_splitterG23ton56n390_splitterG23ton389n390_9_( clk_7 , buf_splitterG23ton56n390_splitterG23ton389n390_10 , 0 , buf_splitterG23ton56n390_splitterG23ton389n390_9 );
buf_AQFP buf_splitterG23ton56n390_splitterG23ton389n390_8_( clk_1 , buf_splitterG23ton56n390_splitterG23ton389n390_9 , 0 , buf_splitterG23ton56n390_splitterG23ton389n390_8 );
buf_AQFP buf_splitterG23ton56n390_splitterG23ton389n390_7_( clk_3 , buf_splitterG23ton56n390_splitterG23ton389n390_8 , 0 , buf_splitterG23ton56n390_splitterG23ton389n390_7 );
buf_AQFP buf_splitterG23ton56n390_splitterG23ton389n390_6_( clk_5 , buf_splitterG23ton56n390_splitterG23ton389n390_7 , 0 , buf_splitterG23ton56n390_splitterG23ton389n390_6 );
buf_AQFP buf_splitterG23ton56n390_splitterG23ton389n390_5_( clk_7 , buf_splitterG23ton56n390_splitterG23ton389n390_6 , 0 , buf_splitterG23ton56n390_splitterG23ton389n390_5 );
buf_AQFP buf_splitterG23ton56n390_splitterG23ton389n390_4_( clk_1 , buf_splitterG23ton56n390_splitterG23ton389n390_5 , 0 , buf_splitterG23ton56n390_splitterG23ton389n390_4 );
buf_AQFP buf_splitterG23ton56n390_splitterG23ton389n390_3_( clk_3 , buf_splitterG23ton56n390_splitterG23ton389n390_4 , 0 , buf_splitterG23ton56n390_splitterG23ton389n390_3 );
buf_AQFP buf_splitterG23ton56n390_splitterG23ton389n390_2_( clk_5 , buf_splitterG23ton56n390_splitterG23ton389n390_3 , 0 , buf_splitterG23ton56n390_splitterG23ton389n390_2 );
buf_AQFP buf_splitterG23ton56n390_splitterG23ton389n390_1_( clk_7 , buf_splitterG23ton56n390_splitterG23ton389n390_2 , 0 , buf_splitterG23ton56n390_splitterG23ton389n390_1 );
buf_AQFP buf_splitterG24ton59n394_splitterG24ton393n394_10_( clk_5 , splitterG24ton59n394 , 0 , buf_splitterG24ton59n394_splitterG24ton393n394_10 );
buf_AQFP buf_splitterG24ton59n394_splitterG24ton393n394_9_( clk_7 , buf_splitterG24ton59n394_splitterG24ton393n394_10 , 0 , buf_splitterG24ton59n394_splitterG24ton393n394_9 );
buf_AQFP buf_splitterG24ton59n394_splitterG24ton393n394_8_( clk_1 , buf_splitterG24ton59n394_splitterG24ton393n394_9 , 0 , buf_splitterG24ton59n394_splitterG24ton393n394_8 );
buf_AQFP buf_splitterG24ton59n394_splitterG24ton393n394_7_( clk_3 , buf_splitterG24ton59n394_splitterG24ton393n394_8 , 0 , buf_splitterG24ton59n394_splitterG24ton393n394_7 );
buf_AQFP buf_splitterG24ton59n394_splitterG24ton393n394_6_( clk_5 , buf_splitterG24ton59n394_splitterG24ton393n394_7 , 0 , buf_splitterG24ton59n394_splitterG24ton393n394_6 );
buf_AQFP buf_splitterG24ton59n394_splitterG24ton393n394_5_( clk_7 , buf_splitterG24ton59n394_splitterG24ton393n394_6 , 0 , buf_splitterG24ton59n394_splitterG24ton393n394_5 );
buf_AQFP buf_splitterG24ton59n394_splitterG24ton393n394_4_( clk_1 , buf_splitterG24ton59n394_splitterG24ton393n394_5 , 0 , buf_splitterG24ton59n394_splitterG24ton393n394_4 );
buf_AQFP buf_splitterG24ton59n394_splitterG24ton393n394_3_( clk_3 , buf_splitterG24ton59n394_splitterG24ton393n394_4 , 0 , buf_splitterG24ton59n394_splitterG24ton393n394_3 );
buf_AQFP buf_splitterG24ton59n394_splitterG24ton393n394_2_( clk_5 , buf_splitterG24ton59n394_splitterG24ton393n394_3 , 0 , buf_splitterG24ton59n394_splitterG24ton393n394_2 );
buf_AQFP buf_splitterG24ton59n394_splitterG24ton393n394_1_( clk_7 , buf_splitterG24ton59n394_splitterG24ton393n394_2 , 0 , buf_splitterG24ton59n394_splitterG24ton393n394_1 );
buf_AQFP buf_splitterG25ton207n399_splitterG25ton398n399_11_( clk_5 , splitterG25ton207n399 , 0 , buf_splitterG25ton207n399_splitterG25ton398n399_11 );
buf_AQFP buf_splitterG25ton207n399_splitterG25ton398n399_10_( clk_7 , buf_splitterG25ton207n399_splitterG25ton398n399_11 , 0 , buf_splitterG25ton207n399_splitterG25ton398n399_10 );
buf_AQFP buf_splitterG25ton207n399_splitterG25ton398n399_9_( clk_1 , buf_splitterG25ton207n399_splitterG25ton398n399_10 , 0 , buf_splitterG25ton207n399_splitterG25ton398n399_9 );
buf_AQFP buf_splitterG25ton207n399_splitterG25ton398n399_8_( clk_3 , buf_splitterG25ton207n399_splitterG25ton398n399_9 , 0 , buf_splitterG25ton207n399_splitterG25ton398n399_8 );
buf_AQFP buf_splitterG25ton207n399_splitterG25ton398n399_7_( clk_5 , buf_splitterG25ton207n399_splitterG25ton398n399_8 , 0 , buf_splitterG25ton207n399_splitterG25ton398n399_7 );
buf_AQFP buf_splitterG25ton207n399_splitterG25ton398n399_6_( clk_7 , buf_splitterG25ton207n399_splitterG25ton398n399_7 , 0 , buf_splitterG25ton207n399_splitterG25ton398n399_6 );
buf_AQFP buf_splitterG25ton207n399_splitterG25ton398n399_5_( clk_1 , buf_splitterG25ton207n399_splitterG25ton398n399_6 , 0 , buf_splitterG25ton207n399_splitterG25ton398n399_5 );
buf_AQFP buf_splitterG25ton207n399_splitterG25ton398n399_4_( clk_3 , buf_splitterG25ton207n399_splitterG25ton398n399_5 , 0 , buf_splitterG25ton207n399_splitterG25ton398n399_4 );
buf_AQFP buf_splitterG25ton207n399_splitterG25ton398n399_3_( clk_5 , buf_splitterG25ton207n399_splitterG25ton398n399_4 , 0 , buf_splitterG25ton207n399_splitterG25ton398n399_3 );
buf_AQFP buf_splitterG25ton207n399_splitterG25ton398n399_2_( clk_7 , buf_splitterG25ton207n399_splitterG25ton398n399_3 , 0 , buf_splitterG25ton207n399_splitterG25ton398n399_2 );
buf_AQFP buf_splitterG25ton207n399_splitterG25ton398n399_1_( clk_1 , buf_splitterG25ton207n399_splitterG25ton398n399_2 , 0 , buf_splitterG25ton207n399_splitterG25ton398n399_1 );
buf_AQFP buf_splitterG26ton210n403_splitterG26ton402n403_11_( clk_5 , splitterG26ton210n403 , 0 , buf_splitterG26ton210n403_splitterG26ton402n403_11 );
buf_AQFP buf_splitterG26ton210n403_splitterG26ton402n403_10_( clk_7 , buf_splitterG26ton210n403_splitterG26ton402n403_11 , 0 , buf_splitterG26ton210n403_splitterG26ton402n403_10 );
buf_AQFP buf_splitterG26ton210n403_splitterG26ton402n403_9_( clk_1 , buf_splitterG26ton210n403_splitterG26ton402n403_10 , 0 , buf_splitterG26ton210n403_splitterG26ton402n403_9 );
buf_AQFP buf_splitterG26ton210n403_splitterG26ton402n403_8_( clk_3 , buf_splitterG26ton210n403_splitterG26ton402n403_9 , 0 , buf_splitterG26ton210n403_splitterG26ton402n403_8 );
buf_AQFP buf_splitterG26ton210n403_splitterG26ton402n403_7_( clk_5 , buf_splitterG26ton210n403_splitterG26ton402n403_8 , 0 , buf_splitterG26ton210n403_splitterG26ton402n403_7 );
buf_AQFP buf_splitterG26ton210n403_splitterG26ton402n403_6_( clk_7 , buf_splitterG26ton210n403_splitterG26ton402n403_7 , 0 , buf_splitterG26ton210n403_splitterG26ton402n403_6 );
buf_AQFP buf_splitterG26ton210n403_splitterG26ton402n403_5_( clk_1 , buf_splitterG26ton210n403_splitterG26ton402n403_6 , 0 , buf_splitterG26ton210n403_splitterG26ton402n403_5 );
buf_AQFP buf_splitterG26ton210n403_splitterG26ton402n403_4_( clk_3 , buf_splitterG26ton210n403_splitterG26ton402n403_5 , 0 , buf_splitterG26ton210n403_splitterG26ton402n403_4 );
buf_AQFP buf_splitterG26ton210n403_splitterG26ton402n403_3_( clk_5 , buf_splitterG26ton210n403_splitterG26ton402n403_4 , 0 , buf_splitterG26ton210n403_splitterG26ton402n403_3 );
buf_AQFP buf_splitterG26ton210n403_splitterG26ton402n403_2_( clk_7 , buf_splitterG26ton210n403_splitterG26ton402n403_3 , 0 , buf_splitterG26ton210n403_splitterG26ton402n403_2 );
buf_AQFP buf_splitterG26ton210n403_splitterG26ton402n403_1_( clk_1 , buf_splitterG26ton210n403_splitterG26ton402n403_2 , 0 , buf_splitterG26ton210n403_splitterG26ton402n403_1 );
buf_AQFP buf_splitterG27ton210n407_splitterG27ton406n407_11_( clk_5 , splitterG27ton210n407 , 0 , buf_splitterG27ton210n407_splitterG27ton406n407_11 );
buf_AQFP buf_splitterG27ton210n407_splitterG27ton406n407_10_( clk_7 , buf_splitterG27ton210n407_splitterG27ton406n407_11 , 0 , buf_splitterG27ton210n407_splitterG27ton406n407_10 );
buf_AQFP buf_splitterG27ton210n407_splitterG27ton406n407_9_( clk_1 , buf_splitterG27ton210n407_splitterG27ton406n407_10 , 0 , buf_splitterG27ton210n407_splitterG27ton406n407_9 );
buf_AQFP buf_splitterG27ton210n407_splitterG27ton406n407_8_( clk_3 , buf_splitterG27ton210n407_splitterG27ton406n407_9 , 0 , buf_splitterG27ton210n407_splitterG27ton406n407_8 );
buf_AQFP buf_splitterG27ton210n407_splitterG27ton406n407_7_( clk_5 , buf_splitterG27ton210n407_splitterG27ton406n407_8 , 0 , buf_splitterG27ton210n407_splitterG27ton406n407_7 );
buf_AQFP buf_splitterG27ton210n407_splitterG27ton406n407_6_( clk_7 , buf_splitterG27ton210n407_splitterG27ton406n407_7 , 0 , buf_splitterG27ton210n407_splitterG27ton406n407_6 );
buf_AQFP buf_splitterG27ton210n407_splitterG27ton406n407_5_( clk_1 , buf_splitterG27ton210n407_splitterG27ton406n407_6 , 0 , buf_splitterG27ton210n407_splitterG27ton406n407_5 );
buf_AQFP buf_splitterG27ton210n407_splitterG27ton406n407_4_( clk_3 , buf_splitterG27ton210n407_splitterG27ton406n407_5 , 0 , buf_splitterG27ton210n407_splitterG27ton406n407_4 );
buf_AQFP buf_splitterG27ton210n407_splitterG27ton406n407_3_( clk_5 , buf_splitterG27ton210n407_splitterG27ton406n407_4 , 0 , buf_splitterG27ton210n407_splitterG27ton406n407_3 );
buf_AQFP buf_splitterG27ton210n407_splitterG27ton406n407_2_( clk_7 , buf_splitterG27ton210n407_splitterG27ton406n407_3 , 0 , buf_splitterG27ton210n407_splitterG27ton406n407_2 );
buf_AQFP buf_splitterG27ton210n407_splitterG27ton406n407_1_( clk_1 , buf_splitterG27ton210n407_splitterG27ton406n407_2 , 0 , buf_splitterG27ton210n407_splitterG27ton406n407_1 );
buf_AQFP buf_splitterG28ton207n411_splitterG28ton410n411_11_( clk_5 , splitterG28ton207n411 , 0 , buf_splitterG28ton207n411_splitterG28ton410n411_11 );
buf_AQFP buf_splitterG28ton207n411_splitterG28ton410n411_10_( clk_7 , buf_splitterG28ton207n411_splitterG28ton410n411_11 , 0 , buf_splitterG28ton207n411_splitterG28ton410n411_10 );
buf_AQFP buf_splitterG28ton207n411_splitterG28ton410n411_9_( clk_1 , buf_splitterG28ton207n411_splitterG28ton410n411_10 , 0 , buf_splitterG28ton207n411_splitterG28ton410n411_9 );
buf_AQFP buf_splitterG28ton207n411_splitterG28ton410n411_8_( clk_3 , buf_splitterG28ton207n411_splitterG28ton410n411_9 , 0 , buf_splitterG28ton207n411_splitterG28ton410n411_8 );
buf_AQFP buf_splitterG28ton207n411_splitterG28ton410n411_7_( clk_5 , buf_splitterG28ton207n411_splitterG28ton410n411_8 , 0 , buf_splitterG28ton207n411_splitterG28ton410n411_7 );
buf_AQFP buf_splitterG28ton207n411_splitterG28ton410n411_6_( clk_7 , buf_splitterG28ton207n411_splitterG28ton410n411_7 , 0 , buf_splitterG28ton207n411_splitterG28ton410n411_6 );
buf_AQFP buf_splitterG28ton207n411_splitterG28ton410n411_5_( clk_1 , buf_splitterG28ton207n411_splitterG28ton410n411_6 , 0 , buf_splitterG28ton207n411_splitterG28ton410n411_5 );
buf_AQFP buf_splitterG28ton207n411_splitterG28ton410n411_4_( clk_3 , buf_splitterG28ton207n411_splitterG28ton410n411_5 , 0 , buf_splitterG28ton207n411_splitterG28ton410n411_4 );
buf_AQFP buf_splitterG28ton207n411_splitterG28ton410n411_3_( clk_5 , buf_splitterG28ton207n411_splitterG28ton410n411_4 , 0 , buf_splitterG28ton207n411_splitterG28ton410n411_3 );
buf_AQFP buf_splitterG28ton207n411_splitterG28ton410n411_2_( clk_7 , buf_splitterG28ton207n411_splitterG28ton410n411_3 , 0 , buf_splitterG28ton207n411_splitterG28ton410n411_2 );
buf_AQFP buf_splitterG28ton207n411_splitterG28ton410n411_1_( clk_1 , buf_splitterG28ton207n411_splitterG28ton410n411_2 , 0 , buf_splitterG28ton207n411_splitterG28ton410n411_1 );
buf_AQFP buf_splitterG29ton195n417_splitterG29ton416n417_10_( clk_5 , splitterG29ton195n417 , 0 , buf_splitterG29ton195n417_splitterG29ton416n417_10 );
buf_AQFP buf_splitterG29ton195n417_splitterG29ton416n417_9_( clk_7 , buf_splitterG29ton195n417_splitterG29ton416n417_10 , 0 , buf_splitterG29ton195n417_splitterG29ton416n417_9 );
buf_AQFP buf_splitterG29ton195n417_splitterG29ton416n417_8_( clk_1 , buf_splitterG29ton195n417_splitterG29ton416n417_9 , 0 , buf_splitterG29ton195n417_splitterG29ton416n417_8 );
buf_AQFP buf_splitterG29ton195n417_splitterG29ton416n417_7_( clk_3 , buf_splitterG29ton195n417_splitterG29ton416n417_8 , 0 , buf_splitterG29ton195n417_splitterG29ton416n417_7 );
buf_AQFP buf_splitterG29ton195n417_splitterG29ton416n417_6_( clk_5 , buf_splitterG29ton195n417_splitterG29ton416n417_7 , 0 , buf_splitterG29ton195n417_splitterG29ton416n417_6 );
buf_AQFP buf_splitterG29ton195n417_splitterG29ton416n417_5_( clk_7 , buf_splitterG29ton195n417_splitterG29ton416n417_6 , 0 , buf_splitterG29ton195n417_splitterG29ton416n417_5 );
buf_AQFP buf_splitterG29ton195n417_splitterG29ton416n417_4_( clk_1 , buf_splitterG29ton195n417_splitterG29ton416n417_5 , 0 , buf_splitterG29ton195n417_splitterG29ton416n417_4 );
buf_AQFP buf_splitterG29ton195n417_splitterG29ton416n417_3_( clk_3 , buf_splitterG29ton195n417_splitterG29ton416n417_4 , 0 , buf_splitterG29ton195n417_splitterG29ton416n417_3 );
buf_AQFP buf_splitterG29ton195n417_splitterG29ton416n417_2_( clk_5 , buf_splitterG29ton195n417_splitterG29ton416n417_3 , 0 , buf_splitterG29ton195n417_splitterG29ton416n417_2 );
buf_AQFP buf_splitterG29ton195n417_splitterG29ton416n417_1_( clk_7 , buf_splitterG29ton195n417_splitterG29ton416n417_2 , 0 , buf_splitterG29ton195n417_splitterG29ton416n417_1 );
buf_AQFP buf_splitterG3ton239n292_splitterG3ton291n292_11_( clk_6 , splitterG3ton239n292 , 0 , buf_splitterG3ton239n292_splitterG3ton291n292_11 );
buf_AQFP buf_splitterG3ton239n292_splitterG3ton291n292_10_( clk_8 , buf_splitterG3ton239n292_splitterG3ton291n292_11 , 0 , buf_splitterG3ton239n292_splitterG3ton291n292_10 );
buf_AQFP buf_splitterG3ton239n292_splitterG3ton291n292_9_( clk_2 , buf_splitterG3ton239n292_splitterG3ton291n292_10 , 0 , buf_splitterG3ton239n292_splitterG3ton291n292_9 );
buf_AQFP buf_splitterG3ton239n292_splitterG3ton291n292_8_( clk_4 , buf_splitterG3ton239n292_splitterG3ton291n292_9 , 0 , buf_splitterG3ton239n292_splitterG3ton291n292_8 );
buf_AQFP buf_splitterG3ton239n292_splitterG3ton291n292_7_( clk_6 , buf_splitterG3ton239n292_splitterG3ton291n292_8 , 0 , buf_splitterG3ton239n292_splitterG3ton291n292_7 );
buf_AQFP buf_splitterG3ton239n292_splitterG3ton291n292_6_( clk_8 , buf_splitterG3ton239n292_splitterG3ton291n292_7 , 0 , buf_splitterG3ton239n292_splitterG3ton291n292_6 );
buf_AQFP buf_splitterG3ton239n292_splitterG3ton291n292_5_( clk_2 , buf_splitterG3ton239n292_splitterG3ton291n292_6 , 0 , buf_splitterG3ton239n292_splitterG3ton291n292_5 );
buf_AQFP buf_splitterG3ton239n292_splitterG3ton291n292_4_( clk_4 , buf_splitterG3ton239n292_splitterG3ton291n292_5 , 0 , buf_splitterG3ton239n292_splitterG3ton291n292_4 );
buf_AQFP buf_splitterG3ton239n292_splitterG3ton291n292_3_( clk_6 , buf_splitterG3ton239n292_splitterG3ton291n292_4 , 0 , buf_splitterG3ton239n292_splitterG3ton291n292_3 );
buf_AQFP buf_splitterG3ton239n292_splitterG3ton291n292_2_( clk_8 , buf_splitterG3ton239n292_splitterG3ton291n292_3 , 0 , buf_splitterG3ton239n292_splitterG3ton291n292_2 );
buf_AQFP buf_splitterG3ton239n292_splitterG3ton291n292_1_( clk_2 , buf_splitterG3ton239n292_splitterG3ton291n292_2 , 0 , buf_splitterG3ton239n292_splitterG3ton291n292_1 );
buf_AQFP buf_splitterG30ton195n421_splitterG30ton420n421_10_( clk_5 , splitterG30ton195n421 , 0 , buf_splitterG30ton195n421_splitterG30ton420n421_10 );
buf_AQFP buf_splitterG30ton195n421_splitterG30ton420n421_9_( clk_7 , buf_splitterG30ton195n421_splitterG30ton420n421_10 , 0 , buf_splitterG30ton195n421_splitterG30ton420n421_9 );
buf_AQFP buf_splitterG30ton195n421_splitterG30ton420n421_8_( clk_1 , buf_splitterG30ton195n421_splitterG30ton420n421_9 , 0 , buf_splitterG30ton195n421_splitterG30ton420n421_8 );
buf_AQFP buf_splitterG30ton195n421_splitterG30ton420n421_7_( clk_3 , buf_splitterG30ton195n421_splitterG30ton420n421_8 , 0 , buf_splitterG30ton195n421_splitterG30ton420n421_7 );
buf_AQFP buf_splitterG30ton195n421_splitterG30ton420n421_6_( clk_5 , buf_splitterG30ton195n421_splitterG30ton420n421_7 , 0 , buf_splitterG30ton195n421_splitterG30ton420n421_6 );
buf_AQFP buf_splitterG30ton195n421_splitterG30ton420n421_5_( clk_7 , buf_splitterG30ton195n421_splitterG30ton420n421_6 , 0 , buf_splitterG30ton195n421_splitterG30ton420n421_5 );
buf_AQFP buf_splitterG30ton195n421_splitterG30ton420n421_4_( clk_1 , buf_splitterG30ton195n421_splitterG30ton420n421_5 , 0 , buf_splitterG30ton195n421_splitterG30ton420n421_4 );
buf_AQFP buf_splitterG30ton195n421_splitterG30ton420n421_3_( clk_3 , buf_splitterG30ton195n421_splitterG30ton420n421_4 , 0 , buf_splitterG30ton195n421_splitterG30ton420n421_3 );
buf_AQFP buf_splitterG30ton195n421_splitterG30ton420n421_2_( clk_5 , buf_splitterG30ton195n421_splitterG30ton420n421_3 , 0 , buf_splitterG30ton195n421_splitterG30ton420n421_2 );
buf_AQFP buf_splitterG30ton195n421_splitterG30ton420n421_1_( clk_7 , buf_splitterG30ton195n421_splitterG30ton420n421_2 , 0 , buf_splitterG30ton195n421_splitterG30ton420n421_1 );
buf_AQFP buf_splitterG31ton198n425_splitterG31ton424n425_10_( clk_5 , splitterG31ton198n425 , 0 , buf_splitterG31ton198n425_splitterG31ton424n425_10 );
buf_AQFP buf_splitterG31ton198n425_splitterG31ton424n425_9_( clk_7 , buf_splitterG31ton198n425_splitterG31ton424n425_10 , 0 , buf_splitterG31ton198n425_splitterG31ton424n425_9 );
buf_AQFP buf_splitterG31ton198n425_splitterG31ton424n425_8_( clk_1 , buf_splitterG31ton198n425_splitterG31ton424n425_9 , 0 , buf_splitterG31ton198n425_splitterG31ton424n425_8 );
buf_AQFP buf_splitterG31ton198n425_splitterG31ton424n425_7_( clk_3 , buf_splitterG31ton198n425_splitterG31ton424n425_8 , 0 , buf_splitterG31ton198n425_splitterG31ton424n425_7 );
buf_AQFP buf_splitterG31ton198n425_splitterG31ton424n425_6_( clk_5 , buf_splitterG31ton198n425_splitterG31ton424n425_7 , 0 , buf_splitterG31ton198n425_splitterG31ton424n425_6 );
buf_AQFP buf_splitterG31ton198n425_splitterG31ton424n425_5_( clk_7 , buf_splitterG31ton198n425_splitterG31ton424n425_6 , 0 , buf_splitterG31ton198n425_splitterG31ton424n425_5 );
buf_AQFP buf_splitterG31ton198n425_splitterG31ton424n425_4_( clk_1 , buf_splitterG31ton198n425_splitterG31ton424n425_5 , 0 , buf_splitterG31ton198n425_splitterG31ton424n425_4 );
buf_AQFP buf_splitterG31ton198n425_splitterG31ton424n425_3_( clk_3 , buf_splitterG31ton198n425_splitterG31ton424n425_4 , 0 , buf_splitterG31ton198n425_splitterG31ton424n425_3 );
buf_AQFP buf_splitterG31ton198n425_splitterG31ton424n425_2_( clk_5 , buf_splitterG31ton198n425_splitterG31ton424n425_3 , 0 , buf_splitterG31ton198n425_splitterG31ton424n425_2 );
buf_AQFP buf_splitterG31ton198n425_splitterG31ton424n425_1_( clk_7 , buf_splitterG31ton198n425_splitterG31ton424n425_2 , 0 , buf_splitterG31ton198n425_splitterG31ton424n425_1 );
buf_AQFP buf_splitterG32ton198n429_splitterG32ton428n429_10_( clk_5 , splitterG32ton198n429 , 0 , buf_splitterG32ton198n429_splitterG32ton428n429_10 );
buf_AQFP buf_splitterG32ton198n429_splitterG32ton428n429_9_( clk_7 , buf_splitterG32ton198n429_splitterG32ton428n429_10 , 0 , buf_splitterG32ton198n429_splitterG32ton428n429_9 );
buf_AQFP buf_splitterG32ton198n429_splitterG32ton428n429_8_( clk_1 , buf_splitterG32ton198n429_splitterG32ton428n429_9 , 0 , buf_splitterG32ton198n429_splitterG32ton428n429_8 );
buf_AQFP buf_splitterG32ton198n429_splitterG32ton428n429_7_( clk_3 , buf_splitterG32ton198n429_splitterG32ton428n429_8 , 0 , buf_splitterG32ton198n429_splitterG32ton428n429_7 );
buf_AQFP buf_splitterG32ton198n429_splitterG32ton428n429_6_( clk_5 , buf_splitterG32ton198n429_splitterG32ton428n429_7 , 0 , buf_splitterG32ton198n429_splitterG32ton428n429_6 );
buf_AQFP buf_splitterG32ton198n429_splitterG32ton428n429_5_( clk_7 , buf_splitterG32ton198n429_splitterG32ton428n429_6 , 0 , buf_splitterG32ton198n429_splitterG32ton428n429_5 );
buf_AQFP buf_splitterG32ton198n429_splitterG32ton428n429_4_( clk_1 , buf_splitterG32ton198n429_splitterG32ton428n429_5 , 0 , buf_splitterG32ton198n429_splitterG32ton428n429_4 );
buf_AQFP buf_splitterG32ton198n429_splitterG32ton428n429_3_( clk_3 , buf_splitterG32ton198n429_splitterG32ton428n429_4 , 0 , buf_splitterG32ton198n429_splitterG32ton428n429_3 );
buf_AQFP buf_splitterG32ton198n429_splitterG32ton428n429_2_( clk_5 , buf_splitterG32ton198n429_splitterG32ton428n429_3 , 0 , buf_splitterG32ton198n429_splitterG32ton428n429_2 );
buf_AQFP buf_splitterG32ton198n429_splitterG32ton428n429_1_( clk_7 , buf_splitterG32ton198n429_splitterG32ton428n429_2 , 0 , buf_splitterG32ton198n429_splitterG32ton428n429_1 );
buf_AQFP buf_splitterG4ton80n296_splitterG4ton295n296_12_( clk_5 , splitterG4ton80n296 , 0 , buf_splitterG4ton80n296_splitterG4ton295n296_12 );
buf_AQFP buf_splitterG4ton80n296_splitterG4ton295n296_11_( clk_7 , buf_splitterG4ton80n296_splitterG4ton295n296_12 , 0 , buf_splitterG4ton80n296_splitterG4ton295n296_11 );
buf_AQFP buf_splitterG4ton80n296_splitterG4ton295n296_10_( clk_1 , buf_splitterG4ton80n296_splitterG4ton295n296_11 , 0 , buf_splitterG4ton80n296_splitterG4ton295n296_10 );
buf_AQFP buf_splitterG4ton80n296_splitterG4ton295n296_9_( clk_3 , buf_splitterG4ton80n296_splitterG4ton295n296_10 , 0 , buf_splitterG4ton80n296_splitterG4ton295n296_9 );
buf_AQFP buf_splitterG4ton80n296_splitterG4ton295n296_8_( clk_5 , buf_splitterG4ton80n296_splitterG4ton295n296_9 , 0 , buf_splitterG4ton80n296_splitterG4ton295n296_8 );
buf_AQFP buf_splitterG4ton80n296_splitterG4ton295n296_7_( clk_7 , buf_splitterG4ton80n296_splitterG4ton295n296_8 , 0 , buf_splitterG4ton80n296_splitterG4ton295n296_7 );
buf_AQFP buf_splitterG4ton80n296_splitterG4ton295n296_6_( clk_1 , buf_splitterG4ton80n296_splitterG4ton295n296_7 , 0 , buf_splitterG4ton80n296_splitterG4ton295n296_6 );
buf_AQFP buf_splitterG4ton80n296_splitterG4ton295n296_5_( clk_3 , buf_splitterG4ton80n296_splitterG4ton295n296_6 , 0 , buf_splitterG4ton80n296_splitterG4ton295n296_5 );
buf_AQFP buf_splitterG4ton80n296_splitterG4ton295n296_4_( clk_5 , buf_splitterG4ton80n296_splitterG4ton295n296_5 , 0 , buf_splitterG4ton80n296_splitterG4ton295n296_4 );
buf_AQFP buf_splitterG4ton80n296_splitterG4ton295n296_3_( clk_7 , buf_splitterG4ton80n296_splitterG4ton295n296_4 , 0 , buf_splitterG4ton80n296_splitterG4ton295n296_3 );
buf_AQFP buf_splitterG4ton80n296_splitterG4ton295n296_2_( clk_1 , buf_splitterG4ton80n296_splitterG4ton295n296_3 , 0 , buf_splitterG4ton80n296_splitterG4ton295n296_2 );
buf_AQFP buf_splitterG4ton80n296_splitterG4ton295n296_1_( clk_3 , buf_splitterG4ton80n296_splitterG4ton295n296_2 , 0 , buf_splitterG4ton80n296_splitterG4ton295n296_1 );
buf_AQFP buf_splitterG5ton65n302_splitterG5ton301n302_12_( clk_5 , splitterG5ton65n302 , 0 , buf_splitterG5ton65n302_splitterG5ton301n302_12 );
buf_AQFP buf_splitterG5ton65n302_splitterG5ton301n302_11_( clk_7 , buf_splitterG5ton65n302_splitterG5ton301n302_12 , 0 , buf_splitterG5ton65n302_splitterG5ton301n302_11 );
buf_AQFP buf_splitterG5ton65n302_splitterG5ton301n302_10_( clk_1 , buf_splitterG5ton65n302_splitterG5ton301n302_11 , 0 , buf_splitterG5ton65n302_splitterG5ton301n302_10 );
buf_AQFP buf_splitterG5ton65n302_splitterG5ton301n302_9_( clk_3 , buf_splitterG5ton65n302_splitterG5ton301n302_10 , 0 , buf_splitterG5ton65n302_splitterG5ton301n302_9 );
buf_AQFP buf_splitterG5ton65n302_splitterG5ton301n302_8_( clk_5 , buf_splitterG5ton65n302_splitterG5ton301n302_9 , 0 , buf_splitterG5ton65n302_splitterG5ton301n302_8 );
buf_AQFP buf_splitterG5ton65n302_splitterG5ton301n302_7_( clk_7 , buf_splitterG5ton65n302_splitterG5ton301n302_8 , 0 , buf_splitterG5ton65n302_splitterG5ton301n302_7 );
buf_AQFP buf_splitterG5ton65n302_splitterG5ton301n302_6_( clk_1 , buf_splitterG5ton65n302_splitterG5ton301n302_7 , 0 , buf_splitterG5ton65n302_splitterG5ton301n302_6 );
buf_AQFP buf_splitterG5ton65n302_splitterG5ton301n302_5_( clk_3 , buf_splitterG5ton65n302_splitterG5ton301n302_6 , 0 , buf_splitterG5ton65n302_splitterG5ton301n302_5 );
buf_AQFP buf_splitterG5ton65n302_splitterG5ton301n302_4_( clk_5 , buf_splitterG5ton65n302_splitterG5ton301n302_5 , 0 , buf_splitterG5ton65n302_splitterG5ton301n302_4 );
buf_AQFP buf_splitterG5ton65n302_splitterG5ton301n302_3_( clk_7 , buf_splitterG5ton65n302_splitterG5ton301n302_4 , 0 , buf_splitterG5ton65n302_splitterG5ton301n302_3 );
buf_AQFP buf_splitterG5ton65n302_splitterG5ton301n302_2_( clk_1 , buf_splitterG5ton65n302_splitterG5ton301n302_3 , 0 , buf_splitterG5ton65n302_splitterG5ton301n302_2 );
buf_AQFP buf_splitterG5ton65n302_splitterG5ton301n302_1_( clk_3 , buf_splitterG5ton65n302_splitterG5ton301n302_2 , 0 , buf_splitterG5ton65n302_splitterG5ton301n302_1 );
buf_AQFP buf_splitterG6ton219n306_splitterG6ton305n306_12_( clk_5 , splitterG6ton219n306 , 0 , buf_splitterG6ton219n306_splitterG6ton305n306_12 );
buf_AQFP buf_splitterG6ton219n306_splitterG6ton305n306_11_( clk_7 , buf_splitterG6ton219n306_splitterG6ton305n306_12 , 0 , buf_splitterG6ton219n306_splitterG6ton305n306_11 );
buf_AQFP buf_splitterG6ton219n306_splitterG6ton305n306_10_( clk_1 , buf_splitterG6ton219n306_splitterG6ton305n306_11 , 0 , buf_splitterG6ton219n306_splitterG6ton305n306_10 );
buf_AQFP buf_splitterG6ton219n306_splitterG6ton305n306_9_( clk_3 , buf_splitterG6ton219n306_splitterG6ton305n306_10 , 0 , buf_splitterG6ton219n306_splitterG6ton305n306_9 );
buf_AQFP buf_splitterG6ton219n306_splitterG6ton305n306_8_( clk_5 , buf_splitterG6ton219n306_splitterG6ton305n306_9 , 0 , buf_splitterG6ton219n306_splitterG6ton305n306_8 );
buf_AQFP buf_splitterG6ton219n306_splitterG6ton305n306_7_( clk_7 , buf_splitterG6ton219n306_splitterG6ton305n306_8 , 0 , buf_splitterG6ton219n306_splitterG6ton305n306_7 );
buf_AQFP buf_splitterG6ton219n306_splitterG6ton305n306_6_( clk_1 , buf_splitterG6ton219n306_splitterG6ton305n306_7 , 0 , buf_splitterG6ton219n306_splitterG6ton305n306_6 );
buf_AQFP buf_splitterG6ton219n306_splitterG6ton305n306_5_( clk_3 , buf_splitterG6ton219n306_splitterG6ton305n306_6 , 0 , buf_splitterG6ton219n306_splitterG6ton305n306_5 );
buf_AQFP buf_splitterG6ton219n306_splitterG6ton305n306_4_( clk_5 , buf_splitterG6ton219n306_splitterG6ton305n306_5 , 0 , buf_splitterG6ton219n306_splitterG6ton305n306_4 );
buf_AQFP buf_splitterG6ton219n306_splitterG6ton305n306_3_( clk_7 , buf_splitterG6ton219n306_splitterG6ton305n306_4 , 0 , buf_splitterG6ton219n306_splitterG6ton305n306_3 );
buf_AQFP buf_splitterG6ton219n306_splitterG6ton305n306_2_( clk_1 , buf_splitterG6ton219n306_splitterG6ton305n306_3 , 0 , buf_splitterG6ton219n306_splitterG6ton305n306_2 );
buf_AQFP buf_splitterG6ton219n306_splitterG6ton305n306_1_( clk_3 , buf_splitterG6ton219n306_splitterG6ton305n306_2 , 0 , buf_splitterG6ton219n306_splitterG6ton305n306_1 );
buf_AQFP buf_splitterG7ton239n310_splitterG7ton309n310_11_( clk_6 , splitterG7ton239n310 , 0 , buf_splitterG7ton239n310_splitterG7ton309n310_11 );
buf_AQFP buf_splitterG7ton239n310_splitterG7ton309n310_10_( clk_8 , buf_splitterG7ton239n310_splitterG7ton309n310_11 , 0 , buf_splitterG7ton239n310_splitterG7ton309n310_10 );
buf_AQFP buf_splitterG7ton239n310_splitterG7ton309n310_9_( clk_2 , buf_splitterG7ton239n310_splitterG7ton309n310_10 , 0 , buf_splitterG7ton239n310_splitterG7ton309n310_9 );
buf_AQFP buf_splitterG7ton239n310_splitterG7ton309n310_8_( clk_4 , buf_splitterG7ton239n310_splitterG7ton309n310_9 , 0 , buf_splitterG7ton239n310_splitterG7ton309n310_8 );
buf_AQFP buf_splitterG7ton239n310_splitterG7ton309n310_7_( clk_6 , buf_splitterG7ton239n310_splitterG7ton309n310_8 , 0 , buf_splitterG7ton239n310_splitterG7ton309n310_7 );
buf_AQFP buf_splitterG7ton239n310_splitterG7ton309n310_6_( clk_8 , buf_splitterG7ton239n310_splitterG7ton309n310_7 , 0 , buf_splitterG7ton239n310_splitterG7ton309n310_6 );
buf_AQFP buf_splitterG7ton239n310_splitterG7ton309n310_5_( clk_2 , buf_splitterG7ton239n310_splitterG7ton309n310_6 , 0 , buf_splitterG7ton239n310_splitterG7ton309n310_5 );
buf_AQFP buf_splitterG7ton239n310_splitterG7ton309n310_4_( clk_4 , buf_splitterG7ton239n310_splitterG7ton309n310_5 , 0 , buf_splitterG7ton239n310_splitterG7ton309n310_4 );
buf_AQFP buf_splitterG7ton239n310_splitterG7ton309n310_3_( clk_6 , buf_splitterG7ton239n310_splitterG7ton309n310_4 , 0 , buf_splitterG7ton239n310_splitterG7ton309n310_3 );
buf_AQFP buf_splitterG7ton239n310_splitterG7ton309n310_2_( clk_8 , buf_splitterG7ton239n310_splitterG7ton309n310_3 , 0 , buf_splitterG7ton239n310_splitterG7ton309n310_2 );
buf_AQFP buf_splitterG7ton239n310_splitterG7ton309n310_1_( clk_2 , buf_splitterG7ton239n310_splitterG7ton309n310_2 , 0 , buf_splitterG7ton239n310_splitterG7ton309n310_1 );
buf_AQFP buf_splitterG8ton262n314_splitterG8ton313n314_11_( clk_6 , splitterG8ton262n314 , 0 , buf_splitterG8ton262n314_splitterG8ton313n314_11 );
buf_AQFP buf_splitterG8ton262n314_splitterG8ton313n314_10_( clk_8 , buf_splitterG8ton262n314_splitterG8ton313n314_11 , 0 , buf_splitterG8ton262n314_splitterG8ton313n314_10 );
buf_AQFP buf_splitterG8ton262n314_splitterG8ton313n314_9_( clk_2 , buf_splitterG8ton262n314_splitterG8ton313n314_10 , 0 , buf_splitterG8ton262n314_splitterG8ton313n314_9 );
buf_AQFP buf_splitterG8ton262n314_splitterG8ton313n314_8_( clk_4 , buf_splitterG8ton262n314_splitterG8ton313n314_9 , 0 , buf_splitterG8ton262n314_splitterG8ton313n314_8 );
buf_AQFP buf_splitterG8ton262n314_splitterG8ton313n314_7_( clk_6 , buf_splitterG8ton262n314_splitterG8ton313n314_8 , 0 , buf_splitterG8ton262n314_splitterG8ton313n314_7 );
buf_AQFP buf_splitterG8ton262n314_splitterG8ton313n314_6_( clk_8 , buf_splitterG8ton262n314_splitterG8ton313n314_7 , 0 , buf_splitterG8ton262n314_splitterG8ton313n314_6 );
buf_AQFP buf_splitterG8ton262n314_splitterG8ton313n314_5_( clk_2 , buf_splitterG8ton262n314_splitterG8ton313n314_6 , 0 , buf_splitterG8ton262n314_splitterG8ton313n314_5 );
buf_AQFP buf_splitterG8ton262n314_splitterG8ton313n314_4_( clk_4 , buf_splitterG8ton262n314_splitterG8ton313n314_5 , 0 , buf_splitterG8ton262n314_splitterG8ton313n314_4 );
buf_AQFP buf_splitterG8ton262n314_splitterG8ton313n314_3_( clk_6 , buf_splitterG8ton262n314_splitterG8ton313n314_4 , 0 , buf_splitterG8ton262n314_splitterG8ton313n314_3 );
buf_AQFP buf_splitterG8ton262n314_splitterG8ton313n314_2_( clk_8 , buf_splitterG8ton262n314_splitterG8ton313n314_3 , 0 , buf_splitterG8ton262n314_splitterG8ton313n314_2 );
buf_AQFP buf_splitterG8ton262n314_splitterG8ton313n314_1_( clk_2 , buf_splitterG8ton262n314_splitterG8ton313n314_2 , 0 , buf_splitterG8ton262n314_splitterG8ton313n314_1 );
buf_AQFP buf_splitterG9ton96n321_splitterG9ton320n321_11_( clk_5 , splitterG9ton96n321 , 0 , buf_splitterG9ton96n321_splitterG9ton320n321_11 );
buf_AQFP buf_splitterG9ton96n321_splitterG9ton320n321_10_( clk_7 , buf_splitterG9ton96n321_splitterG9ton320n321_11 , 0 , buf_splitterG9ton96n321_splitterG9ton320n321_10 );
buf_AQFP buf_splitterG9ton96n321_splitterG9ton320n321_9_( clk_1 , buf_splitterG9ton96n321_splitterG9ton320n321_10 , 0 , buf_splitterG9ton96n321_splitterG9ton320n321_9 );
buf_AQFP buf_splitterG9ton96n321_splitterG9ton320n321_8_( clk_3 , buf_splitterG9ton96n321_splitterG9ton320n321_9 , 0 , buf_splitterG9ton96n321_splitterG9ton320n321_8 );
buf_AQFP buf_splitterG9ton96n321_splitterG9ton320n321_7_( clk_5 , buf_splitterG9ton96n321_splitterG9ton320n321_8 , 0 , buf_splitterG9ton96n321_splitterG9ton320n321_7 );
buf_AQFP buf_splitterG9ton96n321_splitterG9ton320n321_6_( clk_7 , buf_splitterG9ton96n321_splitterG9ton320n321_7 , 0 , buf_splitterG9ton96n321_splitterG9ton320n321_6 );
buf_AQFP buf_splitterG9ton96n321_splitterG9ton320n321_5_( clk_1 , buf_splitterG9ton96n321_splitterG9ton320n321_6 , 0 , buf_splitterG9ton96n321_splitterG9ton320n321_5 );
buf_AQFP buf_splitterG9ton96n321_splitterG9ton320n321_4_( clk_3 , buf_splitterG9ton96n321_splitterG9ton320n321_5 , 0 , buf_splitterG9ton96n321_splitterG9ton320n321_4 );
buf_AQFP buf_splitterG9ton96n321_splitterG9ton320n321_3_( clk_5 , buf_splitterG9ton96n321_splitterG9ton320n321_4 , 0 , buf_splitterG9ton96n321_splitterG9ton320n321_3 );
buf_AQFP buf_splitterG9ton96n321_splitterG9ton320n321_2_( clk_7 , buf_splitterG9ton96n321_splitterG9ton320n321_3 , 0 , buf_splitterG9ton96n321_splitterG9ton320n321_2 );
buf_AQFP buf_splitterG9ton96n321_splitterG9ton320n321_1_( clk_1 , buf_splitterG9ton96n321_splitterG9ton320n321_2 , 0 , buf_splitterG9ton96n321_splitterG9ton320n321_1 );
buf_AQFP buf_splittern78ton230n300_splittern78ton277n300_1_( clk_1 , splittern78ton230n300 , 0 , buf_splittern78ton230n300_splittern78ton277n300_1 );
buf_AQFP buf_splittern78ton277n300_splittern78ton337n300_2_( clk_4 , splittern78ton277n300 , 0 , buf_splittern78ton277n300_splittern78ton337n300_2 );
buf_AQFP buf_splittern78ton277n300_splittern78ton337n300_1_( clk_6 , buf_splittern78ton277n300_splittern78ton337n300_2 , 0 , buf_splittern78ton277n300_splittern78ton337n300_1 );
buf_AQFP buf_splittern115ton354n405_splittern115ton388n405_2_( clk_3 , splittern115ton354n405 , 0 , buf_splittern115ton354n405_splittern115ton388n405_2 );
buf_AQFP buf_splittern115ton354n405_splittern115ton388n405_1_( clk_5 , buf_splittern115ton354n405_splittern115ton388n405_2 , 0 , buf_splittern115ton354n405_splittern115ton388n405_1 );
buf_AQFP buf_splittern152ton354n409_splittern152ton392n409_2_( clk_3 , splittern152ton354n409 , 0 , buf_splittern152ton354n409_splittern152ton392n409_2 );
buf_AQFP buf_splittern152ton354n409_splittern152ton392n409_1_( clk_5 , buf_splittern152ton354n409_splittern152ton392n409_2 , 0 , buf_splittern152ton354n409_splittern152ton392n409_1 );
buf_AQFP buf_splittern153ton356n281_splittern153ton317n281_2_( clk_3 , splittern153ton356n281 , 0 , buf_splittern153ton356n281_splittern153ton317n281_2 );
buf_AQFP buf_splittern153ton356n281_splittern153ton317n281_1_( clk_5 , buf_splittern153ton356n281_splittern153ton317n281_2 , 0 , buf_splittern153ton356n281_splittern153ton317n281_1 );
buf_AQFP buf_splittern153ton317n281_n281_1_( clk_8 , splittern153ton317n281 , 0 , buf_splittern153ton317n281_n281_1 );
buf_AQFP buf_splittern172ton357n397_splittern172ton380n397_2_( clk_3 , splittern172ton357n397 , 0 , buf_splittern172ton357n397_splittern172ton380n397_2 );
buf_AQFP buf_splittern172ton357n397_splittern172ton380n397_1_( clk_5 , buf_splittern172ton357n397_splittern172ton380n397_2 , 0 , buf_splittern172ton357n397_splittern172ton380n397_1 );
buf_AQFP buf_splittern191ton357n401_splittern191ton384n401_2_( clk_3 , splittern191ton357n401 , 0 , buf_splittern191ton357n401_splittern191ton384n401_2 );
buf_AQFP buf_splittern191ton357n401_splittern191ton384n401_1_( clk_5 , buf_splittern191ton357n401_splittern191ton384n401_2 , 0 , buf_splittern191ton357n401_splittern191ton384n401_1 );
buf_AQFP buf_splitterfromn192_n280_3_( clk_3 , splitterfromn192 , 0 , buf_splitterfromn192_n280_3 );
buf_AQFP buf_splitterfromn192_n280_2_( clk_5 , buf_splitterfromn192_n280_3 , 0 , buf_splitterfromn192_n280_2 );
buf_AQFP buf_splitterfromn192_n280_1_( clk_7 , buf_splitterfromn192_n280_2 , 0 , buf_splitterfromn192_n280_1 );
buf_AQFP buf_splittern229ton277n304_splittern229ton341n304_3_( clk_3 , splittern229ton277n304 , 0 , buf_splittern229ton277n304_splittern229ton341n304_3 );
buf_AQFP buf_splittern229ton277n304_splittern229ton341n304_2_( clk_5 , buf_splittern229ton277n304_splittern229ton341n304_3 , 0 , buf_splittern229ton277n304_splittern229ton341n304_2 );
buf_AQFP buf_splittern229ton277n304_splittern229ton341n304_1_( clk_7 , buf_splittern229ton277n304_splittern229ton341n304_2 , 0 , buf_splittern229ton277n304_splittern229ton341n304_1 );
buf_AQFP buf_splitterfromn230_n396_3_( clk_3 , splitterfromn230 , 0 , buf_splitterfromn230_n396_3 );
buf_AQFP buf_splitterfromn230_n396_2_( clk_5 , buf_splitterfromn230_n396_3 , 0 , buf_splitterfromn230_n396_2 );
buf_AQFP buf_splitterfromn230_n396_1_( clk_7 , buf_splitterfromn230_n396_2 , 0 , buf_splitterfromn230_n396_1 );
buf_AQFP buf_splittern249ton275n308_splittern249ton345n308_2_( clk_4 , splittern249ton275n308 , 0 , buf_splittern249ton275n308_splittern249ton345n308_2 );
buf_AQFP buf_splittern249ton275n308_splittern249ton345n308_1_( clk_6 , buf_splittern249ton275n308_splittern249ton345n308_2 , 0 , buf_splittern249ton275n308_splittern249ton345n308_1 );
buf_AQFP buf_splitterfromn251_n361_3_( clk_3 , splitterfromn251 , 0 , buf_splitterfromn251_n361_3 );
buf_AQFP buf_splitterfromn251_n361_2_( clk_5 , buf_splitterfromn251_n361_3 , 0 , buf_splitterfromn251_n361_2 );
buf_AQFP buf_splitterfromn251_n361_1_( clk_7 , buf_splitterfromn251_n361_2 , 0 , buf_splitterfromn251_n361_1 );
buf_AQFP buf_splittern272ton273n312_splittern272ton349n312_1_( clk_6 , splittern272ton273n312 , 0 , buf_splittern272ton273n312_splittern272ton349n312_1 );
buf_AQFP buf_splitterfromn274_n360_1_( clk_5 , splitterfromn274 , 0 , buf_splitterfromn274_n360_1 );
buf_AQFP buf_splittern298ton356n299_splittern298ton335n299_1_( clk_3 , splittern298ton356n299 , 0 , buf_splittern298ton356n299_splittern298ton335n299_1 );
buf_AQFP buf_splittern298ton335n299_n299_2_( clk_6 , splittern298ton335n299 , 0 , buf_splittern298ton335n299_n299_2 );
buf_AQFP buf_splittern298ton335n299_n299_1_( clk_8 , buf_splittern298ton335n299_n299_2 , 0 , buf_splittern298ton335n299_n299_1 );
buf_AQFP buf_splittern316ton353n318_splittern316ton335n318_1_( clk_3 , splittern316ton353n318 , 0 , buf_splittern316ton353n318_splittern316ton335n318_1 );
buf_AQFP buf_splittern316ton335n318_n318_1_( clk_7 , splittern316ton335n318 , 0 , buf_splittern316ton335n318_n318_1 );
splitter_AQFP splitterG1ton67n284_( clk_2 , G1 , 0 , splitterG1ton67n284 );
splitter_AQFP splitterG1ton83n284_( clk_3 , splitterG1ton67n284 , 0 , splitterG1ton83n284 );
splitter_AQFP splitterG1ton283n284_( clk_4 , buf_splitterG1ton83n284_splitterG1ton283n284_1 , 0 , splitterG1ton283n284 );
splitter_AQFP splitterG10ton218n325_( clk_2 , G10 , 0 , splitterG10ton218n325 );
splitter_AQFP splitterG10ton219n325_( clk_3 , splitterG10ton218n325 , 0 , splitterG10ton219n325 );
splitter_AQFP splitterG10ton324n325_( clk_3 , buf_splitterG10ton219n325_splitterG10ton324n325_1 , 0 , splitterG10ton324n325 );
splitter_AQFP splitterG11ton95n329_( clk_2 , G11 , 0 , splitterG11ton95n329 );
splitter_AQFP splitterG11ton235n329_( clk_3 , splitterG11ton95n329 , 0 , splitterG11ton235n329 );
splitter_AQFP splitterG11ton328n329_( clk_3 , buf_splitterG11ton235n329_splitterG11ton328n329_1 , 0 , splitterG11ton328n329 );
splitter_AQFP splitterG12ton258n333_( clk_2 , G12 , 0 , splitterG12ton258n333 );
splitter_AQFP splitterG12ton93n333_( clk_3 , splitterG12ton258n333 , 0 , splitterG12ton93n333 );
splitter_AQFP splitterG12ton332n333_( clk_3 , buf_splitterG12ton93n333_splitterG12ton332n333_1 , 0 , splitterG12ton332n333 );
splitter_AQFP splitterG13ton132n339_( clk_2 , G13 , 0 , splitterG13ton132n339 );
splitter_AQFP splitterG13ton65n339_( clk_3 , splitterG13ton132n339 , 0 , splitterG13ton65n339 );
splitter_AQFP splitterG13ton338n339_( clk_2 , buf_splitterG13ton65n339_splitterG13ton338n339_1 , 0 , splitterG13ton338n339 );
splitter_AQFP splitterG14ton129n343_( clk_2 , G14 , 0 , splitterG14ton129n343 );
splitter_AQFP splitterG14ton216n343_( clk_3 , splitterG14ton129n343 , 0 , splitterG14ton216n343 );
splitter_AQFP splitterG14ton342n343_( clk_2 , buf_splitterG14ton216n343_splitterG14ton342n343_1 , 0 , splitterG14ton342n343 );
splitter_AQFP splitterG15ton132n347_( clk_2 , G15 , 0 , splitterG15ton132n347 );
splitter_AQFP splitterG15ton236n347_( clk_4 , splitterG15ton132n347 , 0 , splitterG15ton236n347 );
splitter_AQFP splitterG15ton346n347_( clk_2 , buf_splitterG15ton236n347_splitterG15ton346n347_1 , 0 , splitterG15ton346n347 );
splitter_AQFP splitterG16ton129n351_( clk_2 , G16 , 0 , splitterG16ton129n351 );
splitter_AQFP splitterG16ton262n351_( clk_4 , splitterG16ton129n351 , 0 , splitterG16ton262n351 );
splitter_AQFP splitterG16ton350n351_( clk_2 , buf_splitterG16ton262n351_splitterG16ton350n351_1 , 0 , splitterG16ton350n351 );
splitter_AQFP splitterG17ton161n364_( clk_2 , G17 , 0 , splitterG17ton161n364 );
splitter_AQFP splitterG17ton44n364_( clk_3 , splitterG17ton161n364 , 0 , splitterG17ton44n364 );
splitter_AQFP splitterG17ton363n364_( clk_2 , buf_splitterG17ton44n364_splitterG17ton363n364_1 , 0 , splitterG17ton363n364 );
splitter_AQFP splitterG18ton177n368_( clk_2 , G18 , 0 , splitterG18ton177n368 );
splitter_AQFP splitterG18ton47n368_( clk_3 , splitterG18ton177n368 , 0 , splitterG18ton47n368 );
splitter_AQFP splitterG18ton367n368_( clk_2 , buf_splitterG18ton47n368_splitterG18ton367n368_1 , 0 , splitterG18ton367n368 );
splitter_AQFP splitterG19ton101n372_( clk_2 , G19 , 0 , splitterG19ton101n372 );
splitter_AQFP splitterG19ton44n372_( clk_3 , splitterG19ton101n372 , 0 , splitterG19ton44n372 );
splitter_AQFP splitterG19ton371n372_( clk_2 , buf_splitterG19ton44n372_splitterG19ton371n372_1 , 0 , splitterG19ton371n372 );
splitter_AQFP splitterG2ton215n288_( clk_2 , G2 , 0 , splitterG2ton215n288 );
splitter_AQFP splitterG2ton216n288_( clk_3 , splitterG2ton215n288 , 0 , splitterG2ton216n288 );
splitter_AQFP splitterG2ton287n288_( clk_4 , buf_splitterG2ton216n288_splitterG2ton287n288_1 , 0 , splitterG2ton287n288 );
splitter_AQFP splitterG20ton138n376_( clk_2 , G20 , 0 , splitterG20ton138n376 );
splitter_AQFP splitterG20ton47n376_( clk_3 , splitterG20ton138n376 , 0 , splitterG20ton47n376 );
splitter_AQFP splitterG20ton375n376_( clk_2 , buf_splitterG20ton47n376_splitterG20ton375n376_1 , 0 , splitterG20ton375n376 );
splitter_AQFP splitterG21ton158n382_( clk_2 , G21 , 0 , splitterG21ton158n382 );
splitter_AQFP splitterG21ton59n382_( clk_3 , splitterG21ton158n382 , 0 , splitterG21ton59n382 );
splitter_AQFP splitterG21ton381n382_( clk_8 , buf_splitterG21ton59n382_splitterG21ton381n382_1 , 0 , splitterG21ton381n382 );
splitter_AQFP splitterG22ton180n386_( clk_2 , G22 , 0 , splitterG22ton180n386 );
splitter_AQFP splitterG22ton56n386_( clk_3 , splitterG22ton180n386 , 0 , splitterG22ton56n386 );
splitter_AQFP splitterG22ton385n386_( clk_8 , buf_splitterG22ton56n386_splitterG22ton385n386_1 , 0 , splitterG22ton385n386 );
splitter_AQFP splitterG23ton101n390_( clk_2 , G23 , 0 , splitterG23ton101n390 );
splitter_AQFP splitterG23ton56n390_( clk_3 , splitterG23ton101n390 , 0 , splitterG23ton56n390 );
splitter_AQFP splitterG23ton389n390_( clk_8 , buf_splitterG23ton56n390_splitterG23ton389n390_1 , 0 , splitterG23ton389n390 );
splitter_AQFP splitterG24ton138n394_( clk_2 , G24 , 0 , splitterG24ton138n394 );
splitter_AQFP splitterG24ton59n394_( clk_3 , splitterG24ton138n394 , 0 , splitterG24ton59n394 );
splitter_AQFP splitterG24ton393n394_( clk_8 , buf_splitterG24ton59n394_splitterG24ton393n394_1 , 0 , splitterG24ton393n394 );
splitter_AQFP splitterG25ton158n399_( clk_2 , G25 , 0 , splitterG25ton158n399 );
splitter_AQFP splitterG25ton207n399_( clk_3 , splitterG25ton158n399 , 0 , splitterG25ton207n399 );
splitter_AQFP splitterG25ton398n399_( clk_2 , buf_splitterG25ton207n399_splitterG25ton398n399_1 , 0 , splitterG25ton398n399 );
splitter_AQFP splitterG26ton177n403_( clk_2 , G26 , 0 , splitterG26ton177n403 );
splitter_AQFP splitterG26ton210n403_( clk_3 , splitterG26ton177n403 , 0 , splitterG26ton210n403 );
splitter_AQFP splitterG26ton402n403_( clk_2 , buf_splitterG26ton210n403_splitterG26ton402n403_1 , 0 , splitterG26ton402n403 );
splitter_AQFP splitterG27ton104n407_( clk_2 , G27 , 0 , splitterG27ton104n407 );
splitter_AQFP splitterG27ton210n407_( clk_3 , splitterG27ton104n407 , 0 , splitterG27ton210n407 );
splitter_AQFP splitterG27ton406n407_( clk_2 , buf_splitterG27ton210n407_splitterG27ton406n407_1 , 0 , splitterG27ton406n407 );
splitter_AQFP splitterG28ton141n411_( clk_2 , G28 , 0 , splitterG28ton141n411 );
splitter_AQFP splitterG28ton207n411_( clk_3 , splitterG28ton141n411 , 0 , splitterG28ton207n411 );
splitter_AQFP splitterG28ton410n411_( clk_2 , buf_splitterG28ton207n411_splitterG28ton410n411_1 , 0 , splitterG28ton410n411 );
splitter_AQFP splitterG29ton161n417_( clk_2 , G29 , 0 , splitterG29ton161n417 );
splitter_AQFP splitterG29ton195n417_( clk_3 , splitterG29ton161n417 , 0 , splitterG29ton195n417 );
splitter_AQFP splitterG29ton416n417_( clk_8 , buf_splitterG29ton195n417_splitterG29ton416n417_1 , 0 , splitterG29ton416n417 );
splitter_AQFP splitterG3ton79n292_( clk_2 , G3 , 0 , splitterG3ton79n292 );
splitter_AQFP splitterG3ton239n292_( clk_4 , splitterG3ton79n292 , 0 , splitterG3ton239n292 );
splitter_AQFP splitterG3ton291n292_( clk_4 , buf_splitterG3ton239n292_splitterG3ton291n292_1 , 0 , splitterG3ton291n292 );
splitter_AQFP splitterG30ton180n421_( clk_2 , G30 , 0 , splitterG30ton180n421 );
splitter_AQFP splitterG30ton195n421_( clk_3 , splitterG30ton180n421 , 0 , splitterG30ton195n421 );
splitter_AQFP splitterG30ton420n421_( clk_8 , buf_splitterG30ton195n421_splitterG30ton420n421_1 , 0 , splitterG30ton420n421 );
splitter_AQFP splitterG31ton104n425_( clk_2 , G31 , 0 , splitterG31ton104n425 );
splitter_AQFP splitterG31ton198n425_( clk_3 , splitterG31ton104n425 , 0 , splitterG31ton198n425 );
splitter_AQFP splitterG31ton424n425_( clk_8 , buf_splitterG31ton198n425_splitterG31ton424n425_1 , 0 , splitterG31ton424n425 );
splitter_AQFP splitterG32ton141n429_( clk_2 , G32 , 0 , splitterG32ton141n429 );
splitter_AQFP splitterG32ton198n429_( clk_3 , splitterG32ton141n429 , 0 , splitterG32ton198n429 );
splitter_AQFP splitterG32ton428n429_( clk_8 , buf_splitterG32ton198n429_splitterG32ton428n429_1 , 0 , splitterG32ton428n429 );
splitter_AQFP splitterG4ton258n296_( clk_2 , G4 , 0 , splitterG4ton258n296 );
splitter_AQFP splitterG4ton80n296_( clk_3 , splitterG4ton258n296 , 0 , splitterG4ton80n296 );
splitter_AQFP splitterG4ton295n296_( clk_4 , buf_splitterG4ton80n296_splitterG4ton295n296_1 , 0 , splitterG4ton295n296 );
splitter_AQFP splitterG41ton173n231_( clk_2 , G41 , 0 , splitterG41ton173n231 );
splitter_AQFP splitterG41ton125n231_( clk_3 , splitterG41ton173n231 , 0 , splitterG41ton125n231 );
splitter_AQFP splitterG41ton254n231_( clk_4 , splitterG41ton125n231 , 0 , splitterG41ton254n231 );
splitter_AQFP splitterG5ton119n302_( clk_2 , G5 , 0 , splitterG5ton119n302 );
splitter_AQFP splitterG5ton65n302_( clk_3 , splitterG5ton119n302 , 0 , splitterG5ton65n302 );
splitter_AQFP splitterG5ton301n302_( clk_4 , buf_splitterG5ton65n302_splitterG5ton301n302_1 , 0 , splitterG5ton301n302 );
splitter_AQFP splitterG6ton119n306_( clk_2 , G6 , 0 , splitterG6ton119n306 );
splitter_AQFP splitterG6ton219n306_( clk_3 , splitterG6ton119n306 , 0 , splitterG6ton219n306 );
splitter_AQFP splitterG6ton305n306_( clk_4 , buf_splitterG6ton219n306_splitterG6ton305n306_1 , 0 , splitterG6ton305n306 );
splitter_AQFP splitterG7ton116n310_( clk_2 , G7 , 0 , splitterG7ton116n310 );
splitter_AQFP splitterG7ton239n310_( clk_4 , splitterG7ton116n310 , 0 , splitterG7ton239n310 );
splitter_AQFP splitterG7ton309n310_( clk_4 , buf_splitterG7ton239n310_splitterG7ton309n310_1 , 0 , splitterG7ton309n310 );
splitter_AQFP splitterG8ton116n314_( clk_2 , G8 , 0 , splitterG8ton116n314 );
splitter_AQFP splitterG8ton262n314_( clk_4 , splitterG8ton116n314 , 0 , splitterG8ton262n314 );
splitter_AQFP splitterG8ton313n314_( clk_4 , buf_splitterG8ton262n314_splitterG8ton313n314_1 , 0 , splitterG8ton313n314 );
splitter_AQFP splitterG9ton67n321_( clk_2 , G9 , 0 , splitterG9ton67n321 );
splitter_AQFP splitterG9ton96n321_( clk_3 , splitterG9ton67n321 , 0 , splitterG9ton96n321 );
splitter_AQFP splitterG9ton320n321_( clk_3 , buf_splitterG9ton96n321_splitterG9ton320n321_1 , 0 , splitterG9ton320n321 );
splitter_AQFP splitterfromn42_( clk_8 , buf_n42_splitterfromn42_1 , 0 , splitterfromn42 );
splitter_AQFP splitterfromn45_( clk_6 , n45 , 0 , splitterfromn45 );
splitter_AQFP splitterfromn48_( clk_6 , n48 , 0 , splitterfromn48 );
splitter_AQFP splittern51ton232n53_( clk_1 , n51 , 0 , splittern51ton232n53 );
splitter_AQFP splitterfromn54_( clk_4 , n54 , 0 , splitterfromn54 );
splitter_AQFP splitterfromn57_( clk_6 , n57 , 0 , splitterfromn57 );
splitter_AQFP splitterfromn60_( clk_6 , n60 , 0 , splitterfromn60 );
splitter_AQFP splittern63ton255n74_( clk_1 , n63 , 0 , splittern63ton255n74 );
splitter_AQFP splitterfromn66_( clk_6 , n66 , 0 , splitterfromn66 );
splitter_AQFP splitterfromn69_( clk_5 , n69 , 0 , splitterfromn69 );
splitter_AQFP splitterfromn72_( clk_1 , n72 , 0 , splitterfromn72 );
splitter_AQFP splitterfromn75_( clk_4 , n75 , 0 , splitterfromn75 );
splitter_AQFP splittern78ton230n300_( clk_7 , n78 , 0 , splittern78ton230n300 );
splitter_AQFP splittern78ton277n300_( clk_2 , buf_splittern78ton230n300_splittern78ton277n300_1 , 0 , splittern78ton277n300 );
splitter_AQFP splittern78ton337n300_( clk_8 , buf_splittern78ton277n300_splittern78ton337n300_1 , 0 , splittern78ton337n300 );
splitter_AQFP splittern78ton319n300_( clk_2 , splittern78ton337n300 , 0 , splittern78ton319n300 );
splitter_AQFP splitterfromn81_( clk_6 , n81 , 0 , splitterfromn81 );
splitter_AQFP splitterfromn84_( clk_6 , n84 , 0 , splitterfromn84 );
splitter_AQFP splittern87ton155n90_( clk_1 , n87 , 0 , splittern87ton155n90 );
splitter_AQFP splitterfromn88_( clk_8 , buf_n88_splitterfromn88_1 , 0 , splitterfromn88 );
splitter_AQFP splitterfromn91_( clk_4 , n91 , 0 , splitterfromn91 );
splitter_AQFP splitterfromn94_( clk_6 , n94 , 0 , splitterfromn94 );
splitter_AQFP splitterfromn97_( clk_6 , n97 , 0 , splitterfromn97 );
splitter_AQFP splittern100ton110n175_( clk_1 , n100 , 0 , splittern100ton110n175 );
splitter_AQFP splitterfromn103_( clk_5 , n103 , 0 , splitterfromn103 );
splitter_AQFP splitterfromn106_( clk_5 , n106 , 0 , splitterfromn106 );
splitter_AQFP splitterfromn109_( clk_8 , n109 , 0 , splitterfromn109 );
splitter_AQFP splitterfromn112_( clk_4 , n112 , 0 , splitterfromn112 );
splitter_AQFP splittern115ton153n405_( clk_7 , n115 , 0 , splittern115ton153n405 );
splitter_AQFP splittern115ton354n405_( clk_1 , splittern115ton153n405 , 0 , splittern115ton354n405 );
splitter_AQFP splittern115ton388n405_( clk_6 , buf_splittern115ton354n405_splittern115ton388n405_1 , 0 , splittern115ton388n405 );
splitter_AQFP splittern115ton370n405_( clk_8 , splittern115ton388n405 , 0 , splittern115ton370n405 );
splitter_AQFP splitterfromn118_( clk_5 , n118 , 0 , splitterfromn118 );
splitter_AQFP splitterfromn121_( clk_5 , n121 , 0 , splitterfromn121 );
splitter_AQFP splittern124ton126n168_( clk_8 , n124 , 0 , splittern124ton126n168 );
splitter_AQFP splitterfromn125_( clk_7 , buf_n125_splitterfromn125_1 , 0 , splitterfromn125 );
splitter_AQFP splitterfromn128_( clk_3 , n128 , 0 , splitterfromn128 );
splitter_AQFP splitterfromn131_( clk_5 , n131 , 0 , splitterfromn131 );
splitter_AQFP splitterfromn134_( clk_5 , n134 , 0 , splitterfromn134 );
splitter_AQFP splittern137ton147n187_( clk_8 , n137 , 0 , splittern137ton147n187 );
splitter_AQFP splitterfromn140_( clk_5 , n140 , 0 , splitterfromn140 );
splitter_AQFP splitterfromn143_( clk_5 , n143 , 0 , splitterfromn143 );
splitter_AQFP splitterfromn146_( clk_8 , n146 , 0 , splitterfromn146 );
splitter_AQFP splitterfromn149_( clk_3 , n149 , 0 , splitterfromn149 );
splitter_AQFP splittern152ton153n409_( clk_7 , n152 , 0 , splittern152ton153n409 );
splitter_AQFP splittern152ton354n409_( clk_1 , splittern152ton153n409 , 0 , splittern152ton354n409 );
splitter_AQFP splittern152ton392n409_( clk_6 , buf_splittern152ton354n409_splittern152ton392n409_1 , 0 , splittern152ton392n409 );
splitter_AQFP splittern152ton374n409_( clk_8 , splittern152ton392n409 , 0 , splittern152ton374n409 );
splitter_AQFP splittern153ton356n281_( clk_1 , n153 , 0 , splittern153ton356n281 );
splitter_AQFP splittern153ton317n281_( clk_6 , buf_splittern153ton356n281_splittern153ton317n281_1 , 0 , splittern153ton317n281 );
splitter_AQFP splitterfromn154_( clk_8 , buf_n154_splitterfromn154_1 , 0 , splitterfromn154 );
splitter_AQFP splitterfromn157_( clk_4 , n157 , 0 , splitterfromn157 );
splitter_AQFP splitterfromn160_( clk_5 , n160 , 0 , splitterfromn160 );
splitter_AQFP splitterfromn163_( clk_5 , n163 , 0 , splitterfromn163 );
splitter_AQFP splitterfromn166_( clk_8 , n166 , 0 , splitterfromn166 );
splitter_AQFP splitterfromn169_( clk_4 , n169 , 0 , splitterfromn169 );
splitter_AQFP splittern172ton192n397_( clk_7 , n172 , 0 , splittern172ton192n397 );
splitter_AQFP splittern172ton357n397_( clk_1 , splittern172ton192n397 , 0 , splittern172ton357n397 );
splitter_AQFP splittern172ton380n397_( clk_6 , buf_splittern172ton357n397_splittern172ton380n397_1 , 0 , splittern172ton380n397 );
splitter_AQFP splittern172ton362n397_( clk_8 , splittern172ton380n397 , 0 , splittern172ton362n397 );
splitter_AQFP splitterfromn173_( clk_8 , buf_n173_splitterfromn173_1 , 0 , splitterfromn173 );
splitter_AQFP splitterfromn176_( clk_4 , n176 , 0 , splitterfromn176 );
splitter_AQFP splitterfromn179_( clk_5 , n179 , 0 , splitterfromn179 );
splitter_AQFP splitterfromn182_( clk_5 , n182 , 0 , splitterfromn182 );
splitter_AQFP splitterfromn185_( clk_8 , n185 , 0 , splitterfromn185 );
splitter_AQFP splitterfromn188_( clk_3 , n188 , 0 , splitterfromn188 );
splitter_AQFP splittern191ton192n401_( clk_7 , n191 , 0 , splittern191ton192n401 );
splitter_AQFP splittern191ton357n401_( clk_1 , splittern191ton192n401 , 0 , splittern191ton357n401 );
splitter_AQFP splittern191ton384n401_( clk_6 , buf_splittern191ton357n401_splittern191ton384n401_1 , 0 , splittern191ton384n401 );
splitter_AQFP splittern191ton366n401_( clk_8 , splittern191ton384n401 , 0 , splittern191ton366n401 );
splitter_AQFP splitterfromn192_( clk_1 , n192 , 0 , splitterfromn192 );
splitter_AQFP splitterfromn193_( clk_8 , buf_n193_splitterfromn193_1 , 0 , splitterfromn193 );
splitter_AQFP splitterfromn196_( clk_6 , n196 , 0 , splitterfromn196 );
splitter_AQFP splitterfromn199_( clk_6 , n199 , 0 , splitterfromn199 );
splitter_AQFP splittern202ton203n268_( clk_1 , n202 , 0 , splittern202ton203n268 );
splitter_AQFP splitterfromn205_( clk_4 , n205 , 0 , splitterfromn205 );
splitter_AQFP splitterfromn208_( clk_6 , n208 , 0 , splitterfromn208 );
splitter_AQFP splitterfromn211_( clk_6 , n211 , 0 , splitterfromn211 );
splitter_AQFP splittern214ton224n245_( clk_1 , n214 , 0 , splittern214ton224n245 );
splitter_AQFP splitterfromn217_( clk_6 , n217 , 0 , splitterfromn217 );
splitter_AQFP splitterfromn220_( clk_6 , n220 , 0 , splitterfromn220 );
splitter_AQFP splitterfromn223_( clk_1 , n223 , 0 , splitterfromn223 );
splitter_AQFP splitterfromn226_( clk_4 , n226 , 0 , splitterfromn226 );
splitter_AQFP splittern229ton230n304_( clk_7 , n229 , 0 , splittern229ton230n304 );
splitter_AQFP splittern229ton277n304_( clk_1 , splittern229ton230n304 , 0 , splittern229ton277n304 );
splitter_AQFP splittern229ton341n304_( clk_8 , buf_splittern229ton277n304_splittern229ton341n304_1 , 0 , splittern229ton341n304 );
splitter_AQFP splittern229ton323n304_( clk_2 , splittern229ton341n304 , 0 , splittern229ton323n304 );
splitter_AQFP splitterfromn230_( clk_1 , n230 , 0 , splitterfromn230 );
splitter_AQFP splitterfromn231_( clk_8 , buf_n231_splitterfromn231_1 , 0 , splitterfromn231 );
splitter_AQFP splitterfromn234_( clk_4 , n234 , 0 , splitterfromn234 );
splitter_AQFP splitterfromn237_( clk_7 , n237 , 0 , splitterfromn237 );
splitter_AQFP splitterfromn240_( clk_7 , n240 , 0 , splitterfromn240 );
splitter_AQFP splitterfromn243_( clk_2 , n243 , 0 , splitterfromn243 );
splitter_AQFP splitterfromn246_( clk_5 , n246 , 0 , splitterfromn246 );
splitter_AQFP splittern249ton250n308_( clk_1 , n249 , 0 , splittern249ton250n308 );
splitter_AQFP splittern249ton275n308_( clk_2 , splittern249ton250n308 , 0 , splittern249ton275n308 );
splitter_AQFP splittern249ton345n308_( clk_8 , buf_splittern249ton275n308_splittern249ton345n308_1 , 0 , splittern249ton345n308 );
splitter_AQFP splittern249ton327n308_( clk_2 , splittern249ton345n308 , 0 , splittern249ton327n308 );
splitter_AQFP splitterfromn250_( clk_3 , n250 , 0 , splitterfromn250 );
splitter_AQFP splitterfromn251_( clk_1 , n251 , 0 , splitterfromn251 );
splitter_AQFP splitterfromn252_( clk_3 , n252 , 0 , splitterfromn252 );
splitter_AQFP splitterfromn254_( clk_8 , buf_n254_splitterfromn254_1 , 0 , splitterfromn254 );
splitter_AQFP splitterfromn257_( clk_4 , n257 , 0 , splitterfromn257 );
splitter_AQFP splitterfromn260_( clk_6 , n260 , 0 , splitterfromn260 );
splitter_AQFP splitterfromn263_( clk_7 , n263 , 0 , splitterfromn263 );
splitter_AQFP splitterfromn266_( clk_2 , n266 , 0 , splitterfromn266 );
splitter_AQFP splitterfromn269_( clk_5 , n269 , 0 , splitterfromn269 );
splitter_AQFP splittern272ton274n312_( clk_8 , n272 , 0 , splittern272ton274n312 );
splitter_AQFP splittern272ton275n312_( clk_2 , splittern272ton274n312 , 0 , splittern272ton275n312 );
splitter_AQFP splittern272ton273n312_( clk_4 , splittern272ton275n312 , 0 , splittern272ton273n312 );
splitter_AQFP splittern272ton349n312_( clk_8 , buf_splittern272ton273n312_splittern272ton349n312_1 , 0 , splittern272ton349n312 );
splitter_AQFP splittern272ton331n312_( clk_2 , splittern272ton349n312 , 0 , splittern272ton331n312 );
splitter_AQFP splitterfromn274_( clk_3 , n274 , 0 , splitterfromn274 );
splitter_AQFP splittern279ton280n336_( clk_7 , n279 , 0 , splittern279ton280n336 );
splitter_AQFP splitterfromn280_( clk_1 , n280 , 0 , splitterfromn280 );
splitter_AQFP splittern281ton282n294_( clk_3 , n281 , 0 , splittern281ton282n294 );
splitter_AQFP splitterfromn282_( clk_5 , n282 , 0 , splitterfromn282 );
splitter_AQFP splitterfromn286_( clk_5 , n286 , 0 , splitterfromn286 );
splitter_AQFP splitterfromn290_( clk_5 , n290 , 0 , splitterfromn290 );
splitter_AQFP splitterfromn294_( clk_5 , n294 , 0 , splitterfromn294 );
splitter_AQFP splittern298ton356n299_( clk_1 , n298 , 0 , splittern298ton356n299 );
splitter_AQFP splittern298ton335n299_( clk_4 , buf_splittern298ton356n299_splittern298ton335n299_1 , 0 , splittern298ton335n299 );
splitter_AQFP splittern299ton300n312_( clk_3 , n299 , 0 , splittern299ton300n312 );
splitter_AQFP splitterfromn300_( clk_5 , n300 , 0 , splitterfromn300 );
splitter_AQFP splitterfromn304_( clk_5 , n304 , 0 , splitterfromn304 );
splitter_AQFP splitterfromn308_( clk_5 , n308 , 0 , splitterfromn308 );
splitter_AQFP splitterfromn312_( clk_5 , n312 , 0 , splitterfromn312 );
splitter_AQFP splittern316ton353n318_( clk_1 , n316 , 0 , splittern316ton353n318 );
splitter_AQFP splittern316ton335n318_( clk_5 , buf_splittern316ton353n318_splittern316ton335n318_1 , 0 , splittern316ton335n318 );
splitter_AQFP splittern318ton319n331_( clk_2 , n318 , 0 , splittern318ton319n331 );
splitter_AQFP splitterfromn319_( clk_4 , n319 , 0 , splitterfromn319 );
splitter_AQFP splitterfromn323_( clk_4 , n323 , 0 , splitterfromn323 );
splitter_AQFP splitterfromn327_( clk_4 , n327 , 0 , splitterfromn327 );
splitter_AQFP splitterfromn331_( clk_4 , n331 , 0 , splitterfromn331 );
splitter_AQFP splittern336ton337n349_( clk_1 , n336 , 0 , splittern336ton337n349 );
splitter_AQFP splitterfromn337_( clk_3 , n337 , 0 , splitterfromn337 );
splitter_AQFP splitterfromn341_( clk_3 , n341 , 0 , splitterfromn341 );
splitter_AQFP splitterfromn345_( clk_3 , n345 , 0 , splitterfromn345 );
splitter_AQFP splitterfromn349_( clk_3 , n349 , 0 , splitterfromn349 );
splitter_AQFP splittern359ton360n414_( clk_5 , n359 , 0 , splittern359ton360n414 );
splitter_AQFP splitterfromn360_( clk_7 , n360 , 0 , splitterfromn360 );
splitter_AQFP splittern361ton362n374_( clk_1 , n361 , 0 , splittern361ton362n374 );
splitter_AQFP splitterfromn362_( clk_3 , n362 , 0 , splitterfromn362 );
splitter_AQFP splitterfromn366_( clk_3 , n366 , 0 , splitterfromn366 );
splitter_AQFP splitterfromn370_( clk_3 , n370 , 0 , splitterfromn370 );
splitter_AQFP splitterfromn374_( clk_3 , n374 , 0 , splitterfromn374 );
splitter_AQFP splittern379ton380n392_( clk_7 , n379 , 0 , splittern379ton380n392 );
splitter_AQFP splitterfromn380_( clk_1 , n380 , 0 , splitterfromn380 );
splitter_AQFP splitterfromn384_( clk_1 , n384 , 0 , splitterfromn384 );
splitter_AQFP splitterfromn388_( clk_1 , n388 , 0 , splitterfromn388 );
splitter_AQFP splitterfromn392_( clk_1 , n392 , 0 , splitterfromn392 );
splitter_AQFP splittern396ton397n409_( clk_1 , n396 , 0 , splittern396ton397n409 );
splitter_AQFP splitterfromn397_( clk_3 , n397 , 0 , splitterfromn397 );
splitter_AQFP splitterfromn401_( clk_3 , n401 , 0 , splitterfromn401 );
splitter_AQFP splitterfromn405_( clk_3 , n405 , 0 , splitterfromn405 );
splitter_AQFP splitterfromn409_( clk_3 , n409 , 0 , splitterfromn409 );
splitter_AQFP splittern414ton415n427_( clk_7 , n414 , 0 , splittern414ton415n427 );
splitter_AQFP splitterfromn415_( clk_1 , n415 , 0 , splitterfromn415 );
splitter_AQFP splitterfromn419_( clk_1 , n419 , 0 , splitterfromn419 );
splitter_AQFP splitterfromn423_( clk_1 , n423 , 0 , splitterfromn423 );
splitter_AQFP splitterfromn427_( clk_1 , n427 , 0 , splitterfromn427 );

endmodule