module top( clk_1 , clk_2 , clk_3 , clk_4 , clk_5 , clk_6 , clk_7 , clk_8 , N1 , N101 , N106 , N111 , N116 , N121 , N126 , N13 , N130 , N135 , N138 , N143 , N146 , N149 , N152 , N153 , N156 , N159 , N165 , N17 , N171 , N177 , N183 , N189 , N195 , N201 , N207 , N210 , N219 , N228 , N237 , N246 , N255 , N259 , N26 , N260 , N261 , N267 , N268 , N29 , N36 , N42 , N51 , N55 , N59 , N68 , N72 , N73 , N74 , N75 , N8 , N80 , N85 , N86 , N87 , N88 , N89 , N90 , N91 , N96 , N388 , N389 , N390 , N391 , N418 , N419 , N420 , N421 , N422 , N423 , N446 , N447 , N448 , N449 , N450 , N767 , N768 , N850 , N863 , N864 , N865 , N866 , N874 , N878 , N879 , N880 );

input N1 , N101 , N106 , N111 , N116 , N121 , N126 , N13 , N130 , N135 , N138 , N143 , N146 , N149 , N152 , N153 , N156 , N159 , N165 , N17 , N171 , N177 , N183 , N189 , N195 , N201 , N207 , N210 , N219 , N228 , N237 , N246 , N255 , N259 , N26 , N260 , N261 , N267 , N268 , N29 , N36 , N42 , N51 , N55 , N59 , N68 , N72 , N73 , N74 , N75 , N8 , N80 , N85 , N86 , N87 , N88 , N89 , N90 , N91 , N96 ;
output N388 , N389 , N390 , N391 , N418 , N419 , N420 , N421 , N422 , N423 , N446 , N447 , N448 , N449 , N450 , N767 , N768 , N850 , N863 , N864 , N865 , N866 , N874 , N878 , N879 , N880 ;
wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , buf_N101_splitterN101ton102n316_1 , buf_N106_splitterN106ton102n289_1 , buf_N111_splitterN111ton105n237_1 , buf_N116_splitterN116ton105n255_1 , buf_N121_splitterN121ton182n97_1 , buf_N121_splitterN121ton182n97_2 , buf_N126_splitterN126ton100n99_1 , buf_N126_splitterN126ton100n99_2 , buf_N13_splitterfromN13_1 , buf_N135_splitterfromN135_1 , buf_N138_splitterN138ton267n291_1 , buf_N138_splitterN138ton267n291_2 , buf_N143_splitterfromN143_1 , buf_N143_splitterfromN143_2 , buf_N143_splitterfromN143_3 , buf_N143_splitterfromN143_4 , buf_N143_splitterfromN143_5 , buf_N146_splitterfromN146_1 , buf_N146_splitterfromN146_2 , buf_N149_splitterfromN149_1 , buf_N149_splitterfromN149_2 , buf_N149_splitterfromN149_3 , buf_N149_splitterfromN149_4 , buf_N152_n291_1 , buf_N152_n291_2 , buf_N152_n291_3 , buf_N153_splitterfromN153_1 , buf_N153_splitterfromN153_2 , buf_N159_splitterN159ton117n330_1 , buf_N165_splitterN165ton129n346_1 , buf_N165_splitterN165ton129n346_2 , buf_N171_splitterN171ton132n361_1 , buf_N171_splitterN171ton132n361_2 , buf_N171_splitterN171ton132n361_3 , buf_N177_splitterN177ton117n315_1 , buf_N177_splitterN177ton117n315_2 , buf_N183_splitterN183ton132n221_1 , buf_N183_splitterN183ton132n221_2 , buf_N183_splitterN183ton132n221_3 , buf_N189_splitterN189ton123n236_1 , buf_N195_splitterN195ton123n253_1 , buf_N195_splitterN195ton123n253_2 , buf_N195_splitterN195ton123n253_3 , buf_N195_splitterN195ton123n253_4 , buf_N201_splitterN201ton129n180_1 , buf_N207_splitterfromN207_1 , buf_N207_splitterfromN207_2 , buf_N207_splitterfromN207_3 , buf_N207_splitterfromN207_4 , buf_N207_splitterfromN207_5 , buf_N207_splitterfromN207_6 , buf_N210_splitterN210ton182n360_1 , buf_N219_splitterN219ton171n355_1 , buf_N219_splitterN219ton171n355_2 , buf_N219_splitterN219ton171n355_3 , buf_N219_splitterN219ton171n355_4 , buf_N219_splitterN219ton171n355_5 , buf_N228_splitterN228ton173n357_1 , buf_N228_splitterN228ton173n357_2 , buf_N228_splitterN228ton173n357_3 , buf_N228_splitterN228ton173n357_4 , buf_N228_splitterN228ton173n357_5 , buf_N228_splitterN228ton173n357_6 , buf_N228_splitterN228ton173n357_7 , buf_N228_splitterN228ton173n357_8 , buf_N237_splitterN237ton174n358_1 , buf_N246_splitterN246ton175n359_1 , buf_N246_splitterN246ton175n359_2 , buf_N246_splitterN246ton175n359_3 , buf_N246_splitterN246ton175n359_4 , buf_N246_splitterN246ton175n359_5 , buf_N255_splitterN255ton181n254_1 , buf_N259_n238_1 , buf_N259_n238_2 , buf_N260_n254_1 , buf_N260_n254_2 , buf_N261_splitterN261ton169n201_1 , buf_N261_splitterN261ton169n201_2 , buf_N261_splitterN261ton169n201_3 , buf_N261_splitterN261ton169n201_4 , buf_N267_n181_1 , buf_N267_n181_2 , buf_N268_splitterN268ton152n331_1 , buf_N51_splitterN51ton159n81_1 , buf_N55_splitterN55ton151n82_1 , buf_N55_splitterN55ton151n82_2 , buf_N72_n176_1 , buf_N72_n176_2 , buf_N73_n177_1 , buf_N73_n177_2 , buf_N74_n87_1 , buf_N74_n87_2 , buf_N74_n87_3 , buf_N80_splitterN80ton149n76_1 , buf_N80_splitterN80ton149n76_2 , buf_N89_n89_1 , buf_N89_n89_2 , buf_N90_n79_1 , buf_N90_n79_2 , buf_N90_n79_3 , buf_N90_n79_4 , buf_N91_splitterN91ton262n94_1 , buf_N91_splitterN91ton262n94_2 , buf_n62_N388_1 , buf_n62_N388_2 , buf_n62_N388_3 , buf_n62_N388_4 , buf_n62_N388_5 , buf_n62_N388_6 , buf_n62_N388_7 , buf_n62_N388_8 , buf_n62_N388_9 , buf_n62_N388_10 , buf_n62_N388_11 , buf_n62_N388_12 , buf_n62_N388_13 , buf_n62_N388_14 , buf_n62_N388_15 , buf_n62_N388_16 , buf_n62_N388_17 , buf_n62_N388_18 , buf_n63_splitterfromn63_1 , buf_n63_splitterfromn63_2 , buf_n64_N389_1 , buf_n64_N389_2 , buf_n64_N389_3 , buf_n64_N389_4 , buf_n64_N389_5 , buf_n64_N389_6 , buf_n64_N389_7 , buf_n64_N389_8 , buf_n64_N389_9 , buf_n64_N389_10 , buf_n64_N389_11 , buf_n64_N389_12 , buf_n64_N389_13 , buf_n64_N389_14 , buf_n64_N389_15 , buf_n64_N389_16 , buf_n64_N389_17 , buf_n64_N389_18 , buf_n65_splittern65toN390n80_1 , buf_n65_splittern65toN390n80_2 , buf_n65_splittern65toN390n80_3 , buf_n65_splittern65toN390n80_4 , buf_n65_splittern65toN390n80_5 , buf_n65_splittern65toN390n80_6 , buf_n65_splittern65toN390n80_7 , buf_n65_splittern65toN390n80_8 , buf_n65_splittern65toN390n80_9 , buf_n65_splittern65toN390n80_10 , buf_n65_splittern65toN390n80_11 , buf_n65_splittern65toN390n80_12 , buf_n65_splittern65toN390n80_13 , buf_n65_splittern65toN390n80_14 , buf_n65_splittern65toN390n80_15 , buf_n66_N391_1 , buf_n66_N391_2 , buf_n66_N391_3 , buf_n66_N391_4 , buf_n66_N391_5 , buf_n66_N391_6 , buf_n66_N391_7 , buf_n66_N391_8 , buf_n66_N391_9 , buf_n66_N391_10 , buf_n66_N391_11 , buf_n66_N391_12 , buf_n66_N391_13 , buf_n66_N391_14 , buf_n66_N391_15 , buf_n66_N391_16 , buf_n66_N391_17 , buf_n66_N391_18 , buf_n66_N391_19 , buf_n66_N391_20 , buf_n66_N391_21 , buf_n67_splittern67ton160n83_1 , buf_n68_splitterfromn68_1 , buf_n68_splitterfromn68_2 , buf_n68_splitterfromn68_3 , buf_n68_splitterfromn68_4 , buf_n69_N418_1 , buf_n69_N418_2 , buf_n69_N418_3 , buf_n69_N418_4 , buf_n69_N418_5 , buf_n69_N418_6 , buf_n69_N418_7 , buf_n71_splitterfromn71_1 , buf_n71_splitterfromn71_2 , buf_n71_splitterfromn71_3 , buf_n71_splitterfromn71_4 , buf_n71_splitterfromn71_5 , buf_n72_N419_1 , buf_n73_splitterfromn73_1 , buf_n74_N420_1 , buf_n74_N420_2 , buf_n74_N420_3 , buf_n74_N420_4 , buf_n74_N420_5 , buf_n74_N420_6 , buf_n74_N420_7 , buf_n74_N420_8 , buf_n74_N420_9 , buf_n74_N420_10 , buf_n74_N420_11 , buf_n74_N420_12 , buf_n74_N420_13 , buf_n74_N420_14 , buf_n74_N420_15 , buf_n74_N420_16 , buf_n74_N420_17 , buf_n74_N420_18 , buf_n76_N421_1 , buf_n76_N421_2 , buf_n76_N421_3 , buf_n76_N421_4 , buf_n76_N421_5 , buf_n76_N421_6 , buf_n76_N421_7 , buf_n76_N421_8 , buf_n76_N421_9 , buf_n77_N422_1 , buf_n77_N422_2 , buf_n77_N422_3 , buf_n77_N422_4 , buf_n77_N422_5 , buf_n77_N422_6 , buf_n77_N422_7 , buf_n77_N422_8 , buf_n77_N422_9 , buf_n77_N422_10 , buf_n77_N422_11 , buf_n77_N422_12 , buf_n77_N422_13 , buf_n77_N422_14 , buf_n77_N422_15 , buf_n77_N422_16 , buf_n77_N422_17 , buf_n77_N422_18 , buf_n77_N422_19 , buf_n77_N422_20 , buf_n77_N422_21 , buf_n77_N422_22 , buf_n77_N422_23 , buf_n77_N422_24 , buf_n79_N423_1 , buf_n79_N423_2 , buf_n79_N423_3 , buf_n79_N423_4 , buf_n79_N423_5 , buf_n79_N423_6 , buf_n79_N423_7 , buf_n79_N423_8 , buf_n79_N423_9 , buf_n79_N423_10 , buf_n79_N423_11 , buf_n79_N423_12 , buf_n79_N423_13 , buf_n79_N423_14 , buf_n79_N423_15 , buf_n79_N423_16 , buf_n79_N423_17 , buf_n79_N423_18 , buf_n79_N423_19 , buf_n79_N423_20 , buf_n79_N423_21 , buf_n80_N446_1 , buf_n84_n85_1 , buf_n84_n85_2 , buf_n84_n85_3 , buf_n84_n85_4 , buf_n84_n85_5 , buf_n84_n85_6 , buf_n84_n85_7 , buf_n84_n85_8 , buf_n84_n85_9 , buf_n84_n85_10 , buf_n84_n85_11 , buf_n84_n85_12 , buf_n84_n85_13 , buf_n84_n85_14 , buf_n84_n85_15 , buf_n84_n85_16 , buf_n85_N448_1 , buf_n85_N448_2 , buf_n85_N448_3 , buf_n87_n88_1 , buf_n88_N449_1 , buf_n88_N449_2 , buf_n88_N449_3 , buf_n88_N449_4 , buf_n88_N449_5 , buf_n88_N449_6 , buf_n88_N449_7 , buf_n88_N449_8 , buf_n88_N449_9 , buf_n88_N449_10 , buf_n88_N449_11 , buf_n88_N449_12 , buf_n88_N449_13 , buf_n88_N449_14 , buf_n88_N449_15 , buf_n88_N449_16 , buf_n88_N449_17 , buf_n89_N450_1 , buf_n89_N450_2 , buf_n89_N450_3 , buf_n89_N450_4 , buf_n89_N450_5 , buf_n89_N450_6 , buf_n89_N450_7 , buf_n89_N450_8 , buf_n89_N450_9 , buf_n89_N450_10 , buf_n89_N450_11 , buf_n89_N450_12 , buf_n89_N450_13 , buf_n89_N450_14 , buf_n89_N450_15 , buf_n89_N450_16 , buf_n89_N450_17 , buf_n89_N450_18 , buf_n89_N450_19 , buf_n89_N450_20 , buf_n89_N450_21 , buf_n89_N450_22 , buf_n89_N450_23 , buf_n89_N450_24 , buf_n89_N450_25 , buf_n89_N450_26 , buf_n89_N450_27 , buf_n89_N450_28 , buf_n89_N450_29 , buf_n89_N450_30 , buf_n89_N450_31 , buf_n89_N450_32 , buf_n89_N450_33 , buf_n89_N450_34 , buf_n89_N450_35 , buf_n89_N450_36 , buf_n93_n95_1 , buf_n94_n95_1 , buf_n95_splitterfromn95_1 , buf_n95_splitterfromn95_2 , buf_n95_splitterfromn95_3 , buf_n113_splitterfromn113_1 , buf_n113_splitterfromn113_2 , buf_n115_n116_1 , buf_n115_n116_2 , buf_n115_n116_3 , buf_n115_n116_4 , buf_n116_N767_1 , buf_n119_splitterfromn119_1 , buf_n122_splitterfromn122_1 , buf_n122_splitterfromn122_2 , buf_n122_splitterfromn122_3 , buf_n140_splitterfromn140_1 , buf_n140_splitterfromn140_2 , buf_n143_N768_1 , buf_n143_N768_2 , buf_n143_N768_3 , buf_n143_N768_4 , buf_n143_N768_5 , buf_n143_N768_6 , buf_n143_N768_7 , buf_n143_N768_8 , buf_n143_N768_9 , buf_n143_N768_10 , buf_n153_n155_1 , buf_n154_n155_1 , buf_n181_n183_1 , buf_n181_n183_2 , buf_n182_n183_1 , buf_n183_n184_1 , buf_n184_n185_1 , buf_n187_n188_1 , buf_n188_N850_1 , buf_n188_N850_2 , buf_n188_N850_3 , buf_n188_N850_4 , buf_n188_N850_5 , buf_n188_N850_6 , buf_n188_N850_7 , buf_n188_N850_8 , buf_n188_N850_9 , buf_n188_N850_10 , buf_n188_N850_11 , buf_n188_N850_12 , buf_n217_n227_1 , buf_n217_n227_2 , buf_n217_n227_3 , buf_n217_n227_4 , buf_n217_n227_5 , buf_n218_n226_1 , buf_n218_n226_2 , buf_n218_n226_3 , buf_n222_n223_1 , buf_n222_n223_2 , buf_n222_n223_3 , buf_n223_n224_1 , buf_n223_n224_2 , buf_n223_n224_3 , buf_n224_n225_1 , buf_n225_n226_1 , buf_n225_n226_2 , buf_n226_n227_1 , buf_n226_n227_2 , buf_n226_n227_3 , buf_n226_n227_4 , buf_n226_n227_5 , buf_n226_n227_6 , buf_n227_N863_1 , buf_n227_N863_2 , buf_n227_N863_3 , buf_n227_N863_4 , buf_n227_N863_5 , buf_n227_N863_6 , buf_n237_n239_1 , buf_n238_n239_1 , buf_n238_n239_2 , buf_n238_n239_3 , buf_n239_n240_1 , buf_n239_n240_2 , buf_n239_n240_3 , buf_n239_n240_4 , buf_n243_n244_1 , buf_n243_n244_2 , buf_n243_n244_3 , buf_n244_N864_1 , buf_n244_N864_2 , buf_n244_N864_3 , buf_n244_N864_4 , buf_n244_N864_5 , buf_n244_N864_6 , buf_n244_N864_7 , buf_n244_N864_8 , buf_n244_N864_9 , buf_n244_N864_10 , buf_n244_N864_11 , buf_n244_N864_12 , buf_n244_N864_13 , buf_n244_N864_14 , buf_n244_N864_15 , buf_n256_n257_1 , buf_n256_n257_2 , buf_n256_n257_3 , buf_n256_n257_4 , buf_n256_n257_5 , buf_n259_n260_1 , buf_n261_N865_1 , buf_n261_N865_2 , buf_n261_N865_3 , buf_n261_N865_4 , buf_n261_N865_5 , buf_n261_N865_6 , buf_n261_N865_7 , buf_n261_N865_8 , buf_n261_N865_9 , buf_n261_N865_10 , buf_n261_N865_11 , buf_n265_n266_1 , buf_n280_splitterfromn280_1 , buf_n280_splitterfromn280_2 , buf_n280_splitterfromn280_3 , buf_n280_splitterfromn280_4 , buf_n306_N866_1 , buf_n306_N866_2 , buf_n307_splitterfromn307_1 , buf_n316_n317_1 , buf_n316_n317_2 , buf_n316_n317_3 , buf_n318_n319_1 , buf_n319_n320_1 , buf_n319_n320_2 , buf_n319_n320_3 , buf_n319_n320_4 , buf_n319_n320_5 , buf_n319_n320_6 , buf_n319_n320_7 , buf_n319_n320_8 , buf_n321_N874_1 , buf_n321_N874_2 , buf_n321_N874_3 , buf_n321_N874_4 , buf_n321_N874_5 , buf_n321_N874_6 , buf_n321_N874_7 , buf_n323_n326_1 , buf_n327_n335_1 , buf_n331_n332_1 , buf_n331_n332_2 , buf_n331_n332_3 , buf_n334_n335_1 , buf_n334_n335_2 , buf_n334_n335_3 , buf_n334_n335_4 , buf_n335_n336_1 , buf_n335_n336_2 , buf_n335_n336_3 , buf_n335_n336_4 , buf_n335_n336_5 , buf_n335_n336_6 , buf_n335_n336_7 , buf_n335_n336_8 , buf_n335_n336_9 , buf_n335_n336_10 , buf_n335_n336_11 , buf_n335_n336_12 , buf_n337_splittern337ton338n342_1 , buf_n337_splittern337ton338n342_2 , buf_n337_splittern337ton338n342_3 , buf_n345_n347_1 , buf_n345_n347_2 , buf_n345_n347_3 , buf_n349_n350_1 , buf_n349_n350_2 , buf_n349_n350_3 , buf_n349_n350_4 , buf_n349_n350_5 , buf_n349_n350_6 , buf_n349_n350_7 , buf_n349_n350_8 , buf_n349_n350_9 , buf_n349_n350_10 , buf_n349_n350_11 , buf_n349_n350_12 , buf_n350_n351_1 , buf_n350_n351_2 , buf_n350_n351_3 , buf_n350_n351_4 , buf_n350_n351_5 , buf_n350_n351_6 , buf_n351_N879_1 , buf_n351_N879_2 , buf_n356_n366_1 , buf_n356_n366_2 , buf_n356_n366_3 , buf_n360_n362_1 , buf_n360_n362_2 , buf_n360_n362_3 , buf_n360_n362_4 , buf_n362_n363_1 , buf_n364_n365_1 , buf_n364_n365_2 , buf_n364_n365_3 , buf_n364_n365_4 , buf_n364_n365_5 , buf_n365_n366_1 , buf_n365_n366_2 , buf_n365_n366_3 , buf_n365_n366_4 , buf_n365_n366_5 , buf_n365_n366_6 , buf_n365_n366_7 , buf_n365_n366_8 , buf_n365_n366_9 , buf_n365_n366_10 , buf_n365_n366_11 , buf_n366_N880_1 , buf_splitterN1ton147n70_n147_1 , buf_splitterN1ton147n70_n147_2 , buf_splitterN1ton147n70_n147_3 , buf_splitterN1ton147n70_n147_4 , buf_splitterN101ton102n316_n281_1 , buf_splitterN101ton102n316_n281_2 , buf_splitterN101ton102n316_n281_3 , buf_splitterN101ton102n316_n316_1 , buf_splitterN106ton102n289_n289_1 , buf_splitterN106ton102n289_n289_2 , buf_splitterN106ton102n289_n289_3 , buf_splitterN111ton105n237_n207_1 , buf_splitterN111ton105n237_n207_2 , buf_splitterN111ton105n237_n207_3 , buf_splitterN116ton105n255_n190_1 , buf_splitterN116ton105n255_n190_2 , buf_splitterN116ton105n255_n255_1 , buf_splitterN121ton182n97_n196_1 , buf_splitterN121ton182n97_n196_2 , buf_splitterN121ton182n97_n196_3 , buf_splitterN126ton100n99_n163_1 , buf_splitterfromN13_n68_1 , buf_splitterN130ton120n91_n120_1 , buf_splitterN130ton120n91_n120_2 , buf_splitterN130ton120n91_n120_3 , buf_splitterN130ton120n91_n120_4 , buf_splitterN130ton120n91_n121_1 , buf_splitterN130ton120n91_n121_2 , buf_splitterN130ton120n91_n121_3 , buf_splitterN130ton120n91_n121_4 , buf_splitterN138ton267n291_n267_1 , buf_splitterN138ton267n291_n283_1 , buf_splitterfromN146_n189_1 , buf_splitterfromN146_n189_2 , buf_splitterfromN146_n274_1 , buf_splitterfromN153_n148_1 , buf_splitterfromN153_n148_2 , buf_splitterfromN153_n290_1 , buf_splitterfromN153_n290_2 , buf_splitterN159ton117n330_n271_1 , buf_splitterN159ton117n330_n271_2 , buf_splitterN159ton117n330_n271_3 , buf_splitterN159ton117n330_n271_4 , buf_splitterN159ton117n330_n271_5 , buf_splitterN165ton129n346_n279_1 , buf_splitterN165ton129n346_n279_2 , buf_splitterN165ton129n346_n279_3 , buf_splitterN165ton129n346_n279_4 , buf_splitterN165ton129n346_n279_5 , buf_splitterN165ton280n346_n280_1 , buf_splitterN17ton146n68_n146_1 , buf_splitterN17ton146n68_n146_2 , buf_splitterN17ton146n68_n146_3 , buf_splitterN17ton159n68_n283_1 , buf_splitterN17ton159n68_n283_2 , buf_splitterN17ton159n68_n283_3 , buf_splitterN17ton159n68_n68_1 , buf_splitterN17ton159n68_n68_2 , buf_splitterN171ton132n361_n287_1 , buf_splitterN171ton132n361_n287_2 , buf_splitterN171ton132n361_n287_3 , buf_splitterN171ton288n361_n288_1 , buf_splitterN177ton117n315_n295_1 , buf_splitterN177ton117n315_n295_2 , buf_splitterN177ton117n315_n295_3 , buf_splitterN177ton117n315_n295_4 , buf_splitterN177ton296n315_n296_1 , buf_splitterN177ton296n315_n296_2 , buf_splitterN183ton132n221_n211_1 , buf_splitterN183ton132n221_n211_2 , buf_splitterN183ton132n221_n211_3 , buf_splitterN183ton212n221_n212_1 , buf_splitterN183ton212n221_n212_2 , buf_splitterN183ton212n221_n212_3 , buf_splitterN189ton123n236_n123_1 , buf_splitterN189ton123n236_n124_1 , buf_splitterN189ton123n236_n124_2 , buf_splitterN189ton123n236_n193_1 , buf_splitterN189ton123n236_n193_2 , buf_splitterN189ton123n236_n193_3 , buf_splitterN189ton123n236_n193_4 , buf_splitterN195ton123n253_n124_1 , buf_splitterN195ton123n253_n199_1 , buf_splitterN195ton123n253_n199_2 , buf_splitterN195ton123n253_n199_3 , buf_splitterN195ton200n253_n200_1 , buf_splitterN195ton200n253_n200_2 , buf_splitterN195ton200n253_n200_3 , buf_splitterN195ton200n253_n253_1 , buf_splitterN201ton129n180_n166_1 , buf_splitterN201ton129n180_n166_2 , buf_splitterN201ton129n180_n166_3 , buf_splitterN201ton129n180_n166_4 , buf_splitterN201ton167n180_n167_1 , buf_splitterN201ton167n180_n167_2 , buf_splitterN201ton167n180_n167_3 , buf_splitterN210ton182n360_n182_1 , buf_splitterN219ton171n355_n171_1 , buf_splitterN219ton171n355_n171_2 , buf_splitterN219ton171n355_n171_3 , buf_splitterN219ton171n355_n217_1 , buf_splitterN219ton171n355_n217_2 , buf_splitterN219ton171n355_n217_3 , buf_splitterN219ton171n355_n217_4 , buf_splitterN219ton171n355_n217_5 , buf_splitterN219ton171n355_n217_6 , buf_splitterN219ton171n355_n217_7 , buf_splitterN219ton232n308_n232_1 , buf_splitterN219ton232n308_n308_1 , buf_splitterN219ton232n308_n308_2 , buf_splitterN219ton232n308_n308_3 , buf_splitterN219ton232n308_n308_4 , buf_splitterN219ton311n355_n325_1 , buf_splitterN219ton311n355_n325_2 , buf_splitterN219ton311n355_n325_3 , buf_splitterN219ton311n355_n325_4 , buf_splitterN219ton311n355_n325_5 , buf_splitterN219ton311n355_n325_6 , buf_splitterN219ton311n355_n340_1 , buf_splitterN219ton311n355_n340_2 , buf_splitterN219ton311n355_n340_3 , buf_splitterN219ton311n355_n340_4 , buf_splitterN219ton311n355_n355_1 , buf_splitterN219ton311n355_n355_2 , buf_splitterN228ton173n357_n173_1 , buf_splitterN228ton173n357_n173_2 , buf_splitterN228ton173n357_n173_3 , buf_splitterN228ton173n357_n218_1 , buf_splitterN228ton173n357_n218_2 , buf_splitterN228ton309n357_n309_1 , buf_splitterN228ton309n357_n309_2 , buf_splitterN228ton309n357_n309_3 , buf_splitterN228ton309n357_n309_4 , buf_splitterN228ton309n357_n309_5 , buf_splitterN228ton309n357_n342_1 , buf_splitterN228ton309n357_n342_2 , buf_splitterN228ton309n357_n342_3 , buf_splitterN228ton309n357_n342_4 , buf_splitterN228ton309n357_n342_5 , buf_splitterN228ton309n357_n342_6 , buf_splitterN228ton309n357_n342_7 , buf_splitterN228ton309n357_n342_8 , buf_splitterN228ton309n357_n342_9 , buf_splitterN228ton309n357_n342_10 , buf_splitterN228ton309n357_n342_11 , buf_splitterN228ton309n357_n357_1 , buf_splitterN237ton174n358_n174_1 , buf_splitterN237ton174n358_n174_2 , buf_splitterN237ton174n358_n174_3 , buf_splitterN237ton174n358_n174_4 , buf_splitterN237ton174n358_n174_5 , buf_splitterN237ton174n358_n219_1 , buf_splitterN237ton174n358_n219_2 , buf_splitterN237ton174n358_n219_3 , buf_splitterN237ton174n358_n219_4 , buf_splitterN237ton174n358_n219_5 , buf_splitterN237ton174n358_n219_6 , buf_splitterN237ton313n358_n313_1 , buf_splitterN237ton313n358_n328_1 , buf_splitterN237ton313n358_n343_1 , buf_splitterN237ton313n358_n358_1 , buf_splitterN237ton313n358_n358_2 , buf_splitterN246ton175n359_n175_1 , buf_splitterN246ton175n359_n220_1 , buf_splitterN261ton169n201_n169_1 , buf_splitterN261ton169n201_n169_2 , buf_splitterN261ton169n201_n169_3 , buf_splitterN261ton169n201_n170_1 , buf_splitterN261ton169n201_n170_2 , buf_splitterN261ton169n201_n170_3 , buf_splitterN261ton169n201_n201_1 , buf_splitterN261ton169n201_n201_2 , buf_splitterN268ton152n331_n152_1 , buf_splitterN268ton152n331_n152_2 , buf_splitterN268ton152n331_n331_1 , buf_splitterN29ton61n84_n84_1 , buf_splitterN42ton153n77_n158_1 , buf_splitterN42ton176n77_n62_1 , buf_splitterN42ton176n77_n65_1 , buf_splitterN42ton176n77_n65_2 , buf_splitterN51ton159n81_n275_1 , buf_splitterN51ton159n81_n275_2 , buf_splitterN55ton151n82_n151_1 , buf_splitterN55ton151n82_n263_1 , buf_splitterN55ton151n82_n263_2 , buf_splitterfromN8_n267_1 , buf_splitterfromN8_n267_2 , buf_splitterfromN8_n267_3 , buf_splitterfromN8_n267_4 , buf_splitterN80ton149n76_n64_1 , buf_splitterN80ton149n76_n64_2 , buf_splitterN80ton149n76_n76_1 , buf_splitterN80ton149n76_n76_2 , buf_splitterN80ton149n76_n76_3 , buf_splitterN80ton149n76_n76_4 , buf_splitterN80ton149n76_n76_5 , buf_splitterN80ton149n76_n76_6 , buf_splitterN80ton149n76_n76_7 , buf_splitterN80ton149n76_n76_8 , buf_splitterN80ton149n76_n76_9 , buf_splitterN80ton149n76_n76_10 , buf_splitterN80ton149n76_n76_11 , buf_splitterN80ton149n76_n76_12 , buf_splitterN91ton262n94_n262_1 , buf_splitterN91ton262n94_n262_2 , buf_splitterN91ton262n94_n345_1 , buf_splitterN91ton262n94_n345_2 , buf_splitterN96ton273n91_n273_1 , buf_splitterN96ton273n91_n273_2 , buf_splitterN96ton273n91_n273_3 , buf_splitterN96ton273n91_n273_4 , buf_splitterN96ton273n91_n273_5 , buf_splitterN96ton273n91_n360_1 , buf_splitterN96ton273n91_n360_2 , buf_splitterfromn61_n62_1 , buf_splitterfromn63_n65_1 , buf_splittern65toN390n80_N390_1 , buf_splittern67ton160n83_n69_1 , buf_splittern67ton160n83_n69_2 , buf_splittern67ton160n83_n69_3 , buf_splittern67ton160n83_n69_4 , buf_splittern67ton160n83_n69_5 , buf_splittern67ton160n83_n69_6 , buf_splittern67ton160n83_n69_7 , buf_splittern67ton160n83_n69_8 , buf_splittern67ton160n83_n69_9 , buf_splittern67ton160n83_n69_10 , buf_splittern67ton160n83_n69_11 , buf_splittern67ton160n83_n83_1 , buf_splitterfromn68_n69_1 , buf_splitterfromn68_n69_2 , buf_splitterfromn68_n69_3 , buf_splitterfromn68_n69_4 , buf_splitterfromn68_n69_5 , buf_splitterfromn68_n69_6 , buf_splitterfromn68_n71_1 , buf_splitterfromn68_n71_2 , buf_splitterfromn68_n71_3 , buf_splitterfromn68_n71_4 , buf_splitterfromn70_n71_1 , buf_splitterfromn70_n71_2 , buf_splitterfromn70_n71_3 , buf_splitterfromn70_n71_4 , buf_splitterfromn70_n71_5 , buf_splitterfromn70_n71_6 , buf_splitterfromn70_n71_7 , buf_splitterfromn70_n71_8 , buf_splitterfromn70_n71_9 , buf_splitterfromn70_n71_10 , buf_splitterfromn70_n71_11 , buf_splitterfromn70_n71_12 , buf_splitterfromn71_n72_1 , buf_splitterfromn71_n80_1 , buf_splitterfromn75_n76_1 , buf_splitterfromn75_n76_2 , buf_splitterfromn75_n76_3 , buf_splitterfromn75_n76_4 , buf_splitterfromn75_n76_5 , buf_splitterfromn75_n76_6 , buf_splitterfromn75_n76_7 , buf_splitterfromn75_n76_8 , buf_splitterfromn75_n76_9 , buf_splitterfromn75_n76_10 , buf_splitterfromn75_n76_11 , buf_splitterfromn75_n76_12 , buf_splitterfromn75_n76_13 , buf_splitterfromn78_n79_1 , buf_splitterfromn78_n79_2 , buf_splitterfromn78_n89_1 , buf_splittern81toN447n156_N447_1 , buf_splittern81toN447n156_N447_2 , buf_splittern81toN447n156_N447_3 , buf_splittern81toN447n156_N447_4 , buf_splittern81toN447n156_N447_5 , buf_splittern81toN447n156_N447_6 , buf_splittern81toN447n156_N447_7 , buf_splittern81toN447n156_N447_8 , buf_splittern81toN447n156_N447_9 , buf_splittern81toN447n156_N447_10 , buf_splittern81toN447n156_N447_11 , buf_splittern81toN447n156_N447_12 , buf_splittern81toN447n156_N447_13 , buf_splittern81toN447n156_N447_14 , buf_splittern81toN447n156_N447_15 , buf_splittern81toN447n156_N447_16 , buf_splittern81toN447n156_N447_17 , buf_splittern81toN447n156_N447_18 , buf_splittern81toN447n156_N447_19 , buf_splittern83ton179n88_n85_1 , buf_splittern83ton179n88_n85_2 , buf_splittern83ton179n88_n85_3 , buf_splittern83ton179n88_n85_4 , buf_splittern83ton179n88_n85_5 , buf_splittern83ton179n88_n85_6 , buf_splittern83ton179n88_n85_7 , buf_splittern83ton179n88_n85_8 , buf_splittern83ton179n88_n85_9 , buf_splittern83ton179n88_n85_10 , buf_splittern83ton179n88_n85_11 , buf_splittern83ton179n88_n85_12 , buf_splittern83ton179n88_n85_13 , buf_splittern83ton179n88_n85_14 , buf_splittern83ton179n88_n85_15 , buf_splittern83ton179n88_n85_16 , buf_splitterfromn95_n114_1 , buf_splitterfromn95_n114_2 , buf_splitterfromn95_n114_3 , buf_splitterfromn95_n114_4 , buf_splitterfromn95_n114_5 , buf_splitterfromn95_n114_6 , buf_splitterfromn95_n114_7 , buf_splitterfromn95_n114_8 , buf_splitterfromn95_n114_9 , buf_splitterfromn95_n114_10 , buf_splitterfromn95_n114_11 , buf_splitterfromn95_n114_12 , buf_splitterfromn95_n115_1 , buf_splitterfromn95_n115_2 , buf_splitterfromn95_n115_3 , buf_splitterfromn95_n115_4 , buf_splitterfromn95_n115_5 , buf_splitterfromn95_n115_6 , buf_splitterfromn95_n115_7 , buf_splitterfromn95_n115_8 , buf_splitterfromn104_n109_1 , buf_splitterfromn113_n114_1 , buf_splitterfromn113_n114_2 , buf_splitterfromn113_n114_3 , buf_splitterfromn113_n114_4 , buf_splitterfromn113_n114_5 , buf_splitterfromn113_n114_6 , buf_splitterfromn113_n114_7 , buf_splitterfromn113_n114_8 , buf_splitterfromn113_n114_9 , buf_splitterfromn113_n114_10 , buf_splitterfromn113_n114_11 , buf_splitterfromn113_n114_12 , buf_splitterfromn113_n114_13 , buf_splitterfromn113_n115_1 , buf_splitterfromn113_n115_2 , buf_splitterfromn113_n115_3 , buf_splitterfromn113_n115_4 , buf_splitterfromn113_n115_5 , buf_splitterfromn122_n141_1 , buf_splitterfromn122_n142_1 , buf_splitterfromn122_n142_2 , buf_splitterfromn122_n142_3 , buf_splitterfromn131_n136_1 , buf_splitterfromn134_n136_1 , buf_splitterfromn144_n145_1 , buf_splitterfromn144_n156_1 , buf_splittern152ton164n210_n210_1 , buf_splittern152ton164n210_n210_2 , buf_splittern193ton206n234_n206_1 , buf_splittern193ton206n234_n206_2 , buf_splittern193ton206n234_n206_3 , buf_splittern193ton206n234_n206_4 , buf_splitterfromn194_n205_1 , buf_splitterfromn194_n205_2 , buf_splitterfromn194_n205_3 , buf_splittern199ton204n251_n204_1 , buf_splitterfromn200_n203_1 , buf_splittern211ton213n298_n298_1 , buf_splittern211ton213n298_n298_2 , buf_splittern211ton213n298_n298_3 , buf_splittern211ton213n298_n298_4 , buf_splitterfromn212_n297_1 , buf_splitterfromn212_n297_2 , buf_splitterfromn212_n297_3 , buf_splitterfromn212_n297_4 , buf_splitterfromn212_n297_5 , buf_splitterfromn212_n297_6 , buf_splittern213ton214n218_n214_1 , buf_splittern213ton214n218_n214_2 , buf_splittern213ton214n218_n214_3 , buf_splittern213ton214n218_n215_1 , buf_splittern213ton214n218_n215_2 , buf_splittern213ton214n218_n215_3 , buf_splittern228ton229n233_n229_1 , buf_splittern228ton229n233_n229_2 , buf_splittern228ton229n233_n230_1 , buf_splittern228ton229n233_n230_2 , buf_splittern271ton306n328_n306_1 , buf_splittern271ton306n328_n306_2 , buf_splittern271ton306n328_n306_3 , buf_splittern271ton306n328_n306_4 , buf_splittern271ton306n328_n306_5 , buf_splittern271ton306n328_n306_6 , buf_splittern271ton306n328_n306_7 , buf_splittern271ton306n328_n306_8 , buf_splittern271ton306n328_n306_9 , buf_splittern271ton306n328_n306_10 , buf_splittern271ton306n328_n306_11 , buf_splittern271ton306n328_n306_12 , buf_splitterfromn272_n305_1 , buf_splitterfromn272_n305_2 , buf_splitterfromn272_n305_3 , buf_splitterfromn272_n305_4 , buf_splitterfromn272_n305_5 , buf_splitterfromn272_n305_6 , buf_splitterfromn272_n305_7 , buf_splitterfromn272_n305_8 , buf_splitterfromn272_n305_9 , buf_splitterfromn272_n305_10 , buf_splittern279ton304n343_n304_1 , buf_splittern279ton304n343_n304_2 , buf_splittern279ton304n343_n304_3 , buf_splittern279ton304n343_n304_4 , buf_splittern279ton304n343_n304_5 , buf_splittern279ton304n343_n304_6 , buf_splittern279ton304n343_n304_7 , buf_splittern279ton304n343_n304_8 , buf_splittern279ton304n343_n304_9 , buf_splittern279ton304n343_n337_1 , buf_splittern279ton304n343_n337_2 , buf_splittern279ton304n343_n337_3 , buf_splitterfromn280_n303_1 , buf_splitterfromn280_n303_2 , buf_splitterfromn280_n303_3 , buf_splitterfromn280_n303_4 , buf_splitterfromn280_n303_5 , buf_splittern287ton302n358_n302_1 , buf_splittern287ton302n358_n302_2 , buf_splittern287ton302n358_n302_3 , buf_splittern287ton302n358_n302_4 , buf_splittern287ton302n358_n302_5 , buf_splittern287ton302n358_n302_6 , buf_splittern287ton302n358_n302_7 , buf_splittern287ton302n358_n302_8 , buf_splittern287ton302n358_n302_9 , buf_splitterfromn288_n301_1 , buf_splitterfromn288_n301_2 , buf_splitterfromn288_n301_3 , buf_splitterfromn288_n301_4 , buf_splitterfromn288_n301_5 , buf_splitterfromn288_n301_6 , buf_splitterfromn288_n301_7 , buf_splitterfromn288_n301_8 , buf_splittern295ton300n313_n300_1 , buf_splittern295ton300n313_n300_2 , buf_splittern295ton300n313_n300_3 , buf_splittern295ton300n313_n300_4 , buf_splittern295ton300n313_n300_5 , buf_splittern295ton300n313_n300_6 , buf_splittern295ton300n313_n307_1 , buf_splitterfromn296_n299_1 , buf_splitterfromn296_n299_2 , buf_splitterfromn296_n299_3 , buf_splitterfromn296_n299_4 , buf_splitterfromn296_n299_5 , buf_splittern298ton299n312_n312_1 , buf_splitterfromn307_n310_1 , buf_splitterfromn307_n310_2 , buf_splitterfromn307_n310_3 , buf_splitterfromn307_n311_1 , buf_splitterfromn307_n311_2 , buf_splittern322ton323n327_n323_1 , buf_splittern322ton323n327_n323_2 , buf_splittern322ton323n327_n323_3 , buf_splittern322ton323n327_n323_4 , buf_splittern322ton323n327_n323_5 , buf_splittern322ton323n327_n323_6 , buf_splittern322ton323n327_n323_7 , buf_splittern322ton323n327_n323_8 , buf_splittern322ton323n327_n323_9 , buf_splittern322ton323n327_n324_1 , buf_splittern322ton323n327_n324_2 , buf_splittern322ton323n327_n324_3 , buf_splittern322ton323n327_n324_4 , buf_splittern322ton323n327_n324_5 , buf_splittern322ton323n327_n324_6 , buf_splittern322ton323n327_n324_7 , buf_splittern322ton323n327_n324_8 , buf_splittern322ton323n327_n324_9 , buf_splittern322ton323n327_n324_10 , buf_splittern337ton338n342_n338_1 , buf_splittern337ton338n342_n338_2 , buf_splittern337ton338n342_n338_3 , buf_splittern337ton338n342_n339_1 , buf_splittern337ton338n342_n339_2 , buf_splittern337ton338n342_n339_3 , buf_splittern337ton338n342_n339_4 , buf_splittern337ton338n342_n339_5 , buf_splittern352ton353n357_n353_1 , buf_splittern352ton353n357_n353_2 , buf_splittern352ton353n357_n353_3 , buf_splittern352ton353n357_n353_4 , buf_splittern352ton353n357_n353_5 , buf_splittern352ton353n357_n353_6 , buf_splittern352ton353n357_n353_7 , buf_splittern352ton353n357_n354_1 , buf_splittern352ton353n357_n354_2 , buf_splittern352ton353n357_n354_3 , buf_splittern352ton353n357_n354_4 , buf_splittern352ton353n357_n354_5 , buf_splittern352ton353n357_n354_6 , splitterN1ton147n70 , splitterN101ton102n316 , splitterN106ton102n289 , splitterN111ton105n237 , splitterN116ton105n255 , splitterN121ton182n97 , splitterN126ton100n99 , splitterfromN13 , splitterN130ton120n91 , splitterfromN135 , splitterN138ton267n291 , splitterfromN143 , splitterfromN146 , splitterfromN149 , splitterfromN153 , splitterN159ton117n330 , splitterN159ton272n330 , splitterN165ton129n346 , splitterN165ton280n346 , splitterN17ton146n68 , splitterN17ton159n68 , splitterN171ton132n361 , splitterN171ton288n361 , splitterN177ton117n315 , splitterN177ton296n315 , splitterN183ton132n221 , splitterN183ton212n221 , splitterN189ton123n236 , splitterN189ton194n236 , splitterN195ton123n253 , splitterN195ton200n253 , splitterN201ton129n180 , splitterN201ton167n180 , splitterfromN207 , splitterN210ton182n360 , splitterN210ton237n255 , splitterN210ton316n360 , splitterN219ton171n355 , splitterN219ton232n308 , splitterN219ton311n355 , splitterN228ton173n357 , splitterN228ton233n250 , splitterN228ton309n357 , splitterN237ton174n358 , splitterN237ton234n251 , splitterN237ton313n358 , splitterN246ton175n359 , splitterN246ton235n252 , splitterN246ton314n359 , splitterN255ton181n254 , splitterN261ton169n201 , splitterN268ton152n331 , splitterN29ton61n84 , splitterfromN36 , splitterN42ton153n77 , splitterN42ton176n77 , splitterN51ton159n81 , splitterN55ton151n82 , splitterN59ton144n86 , splitterfromN68 , splitterfromN75 , splitterfromN8 , splitterN80ton149n76 , splitterN91ton262n94 , splitterN96ton273n91 , splitterfromn61 , splitterfromn63 , splittern65toN390n80 , splittern67ton160n83 , splitterfromn68 , splitterfromn70 , splitterfromn71 , splitterfromn73 , splitterfromn75 , splitterfromn78 , splittern81toN447n156 , splittern83ton179n88 , splitterfromn86 , splitterfromn92 , splitterfromn95 , splitterfromn98 , splitterfromn101 , splitterfromn104 , splitterfromn107 , splitterfromn110 , splitterfromn113 , splitterfromn119 , splitterfromn122 , splitterfromn125 , splitterfromn128 , splitterfromn131 , splitterfromn134 , splitterfromn137 , splitterfromn140 , splitterfromn144 , splitterfromn145 , splittern147ton148n208 , splitterfromn150 , splittern152ton164n210 , splittern162ton163n289 , splittern162ton196n207 , splittern162ton262n289 , splittern165ton166n175 , splitterfromn166 , splittern167ton168n201 , splittern168ton169n173 , splittern179ton180n361 , splittern179ton236n253 , splittern179ton315n361 , splittern192ton193n235 , splittern193ton206n234 , splitterfromn194 , splittern198ton199n252 , splittern199ton204n251 , splitterfromn200 , splittern202ton203n247 , splittern204ton205n230 , splittern206ton214n297 , splittern210ton211n220 , splittern211ton213n298 , splitterfromn212 , splittern213ton214n218 , splittern228ton229n233 , splittern245ton246n250 , splittern263ton264n290 , splittern266ton268n292 , splittern270ton271n329 , splittern271ton306n328 , splitterfromn272 , splittern278ton279n344 , splittern279ton304n343 , splitterfromn280 , splittern286ton287n359 , splittern287ton302n358 , splitterfromn288 , splittern294ton295n314 , splittern295ton300n313 , splitterfromn296 , splittern298ton299n312 , splittern300ton301n354 , splittern302ton303n339 , splittern304ton305n324 , splitterfromn307 , splittern322ton323n327 , splittern337ton338n342 , splittern352ton353n357 ;

PI_AQFP N1_( clk_1 , N1 );
PI_AQFP N101_( clk_1 , N101 );
PI_AQFP N106_( clk_1 , N106 );
PI_AQFP N111_( clk_1 , N111 );
PI_AQFP N116_( clk_1 , N116 );
PI_AQFP N121_( clk_1 , N121 );
PI_AQFP N126_( clk_1 , N126 );
PI_AQFP N13_( clk_1 , N13 );
PI_AQFP N130_( clk_1 , N130 );
PI_AQFP N135_( clk_1 , N135 );
PI_AQFP N138_( clk_1 , N138 );
PI_AQFP N143_( clk_1 , N143 );
PI_AQFP N146_( clk_1 , N146 );
PI_AQFP N149_( clk_1 , N149 );
PI_AQFP N152_( clk_1 , N152 );
PI_AQFP N153_( clk_1 , N153 );
PI_AQFP N156_( clk_1 , N156 );
PI_AQFP N159_( clk_1 , N159 );
PI_AQFP N165_( clk_1 , N165 );
PI_AQFP N17_( clk_1 , N17 );
PI_AQFP N171_( clk_1 , N171 );
PI_AQFP N177_( clk_1 , N177 );
PI_AQFP N183_( clk_1 , N183 );
PI_AQFP N189_( clk_1 , N189 );
PI_AQFP N195_( clk_1 , N195 );
PI_AQFP N201_( clk_1 , N201 );
PI_AQFP N207_( clk_1 , N207 );
PI_AQFP N210_( clk_1 , N210 );
PI_AQFP N219_( clk_1 , N219 );
PI_AQFP N228_( clk_1 , N228 );
PI_AQFP N237_( clk_1 , N237 );
PI_AQFP N246_( clk_1 , N246 );
PI_AQFP N255_( clk_1 , N255 );
PI_AQFP N259_( clk_1 , N259 );
PI_AQFP N26_( clk_1 , N26 );
PI_AQFP N260_( clk_1 , N260 );
PI_AQFP N261_( clk_1 , N261 );
PI_AQFP N267_( clk_1 , N267 );
PI_AQFP N268_( clk_1 , N268 );
PI_AQFP N29_( clk_1 , N29 );
PI_AQFP N36_( clk_1 , N36 );
PI_AQFP N42_( clk_1 , N42 );
PI_AQFP N51_( clk_1 , N51 );
PI_AQFP N55_( clk_1 , N55 );
PI_AQFP N59_( clk_1 , N59 );
PI_AQFP N68_( clk_1 , N68 );
PI_AQFP N72_( clk_1 , N72 );
PI_AQFP N73_( clk_1 , N73 );
PI_AQFP N74_( clk_1 , N74 );
PI_AQFP N75_( clk_1 , N75 );
PI_AQFP N8_( clk_1 , N8 );
PI_AQFP N80_( clk_1 , N80 );
PI_AQFP N85_( clk_1 , N85 );
PI_AQFP N86_( clk_1 , N86 );
PI_AQFP N87_( clk_1 , N87 );
PI_AQFP N88_( clk_1 , N88 );
PI_AQFP N89_( clk_1 , N89 );
PI_AQFP N90_( clk_1 , N90 );
PI_AQFP N91_( clk_1 , N91 );
PI_AQFP N96_( clk_1 , N96 );
and_AQFP n61_( clk_3 , splitterN29ton61n84 , splitterfromN75 , 0 , 0 , n61 );
and_AQFP n62_( clk_1 , buf_splitterN42ton176n77_n62_1 , buf_splitterfromn61_n62_1 , 0 , 0 , n62 );
and_AQFP n63_( clk_3 , splitterN29ton61n84 , splitterfromN36 , 0 , 0 , n63 );
and_AQFP n64_( clk_1 , buf_splitterN80ton149n76_n64_2 , splitterfromn63 , 0 , 0 , n64 );
and_AQFP n65_( clk_3 , buf_splitterN42ton176n77_n65_2 , buf_splitterfromn63_n65_1 , 0 , 0 , n65 );
and_AQFP n66_( clk_3 , N85 , N86 , 0 , 0 , n66 );
and_AQFP n67_( clk_3 , splitterN1ton147n70 , splitterfromN8 , 0 , 0 , n67 );
and_AQFP n68_( clk_7 , buf_splitterfromN13_n68_1 , buf_splitterN17ton159n68_n68_2 , 0 , 0 , n68 );
and_AQFP n69_( clk_5 , buf_splittern67ton160n83_n69_11 , buf_splitterfromn68_n69_6 , 0 , 0 , n69 );
and_AQFP n70_( clk_3 , splitterN1ton147n70 , N26 , 0 , 0 , n70 );
and_AQFP n71_( clk_3 , buf_splitterfromn68_n71_4 , buf_splitterfromn70_n71_12 , 0 , 0 , n71 );
and_AQFP n72_( clk_3 , splittern65toN390n80 , buf_splitterfromn71_n72_1 , 1 , 0 , n72 );
and_AQFP n73_( clk_3 , splitterN59ton144n86 , splitterfromN75 , 0 , 0 , n73 );
and_AQFP n74_( clk_7 , splitterN80ton149n76 , splitterfromn73 , 0 , 0 , n74 );
and_AQFP n75_( clk_3 , splitterfromN36 , splitterN59ton144n86 , 0 , 0 , n75 );
and_AQFP n76_( clk_7 , buf_splitterN80ton149n76_n76_12 , buf_splitterfromn75_n76_13 , 0 , 0 , n76 );
and_AQFP n77_( clk_6 , splitterN42ton176n77 , splitterfromn75 , 0 , 0 , n77 );
or_AQFP n78_( clk_3 , N87 , N88 , 0 , 0 , n78 );
and_AQFP n79_( clk_2 , buf_N90_n79_4 , buf_splitterfromn78_n79_2 , 0 , 0 , n79 );
and_AQFP n80_( clk_3 , splittern65toN390n80 , buf_splitterfromn71_n80_1 , 0 , 0 , n80 );
and_AQFP n81_( clk_5 , splitterN51ton159n81 , splitterfromn70 , 0 , 0 , n81 );
and_AQFP n82_( clk_6 , splitterfromN13 , splitterN55ton151n82 , 0 , 0 , n82 );
and_AQFP n83_( clk_8 , buf_splittern67ton160n83_n83_1 , n82 , 0 , 0 , n83 );
and_AQFP n84_( clk_5 , buf_splitterN29ton61n84_n84_1 , splitterfromN68 , 0 , 0 , n84 );
and_AQFP n85_( clk_6 , buf_splittern83ton179n88_n85_16 , buf_n84_n85_16 , 0 , 0 , n85 );
and_AQFP n86_( clk_4 , splitterN59ton144n86 , splitterfromN68 , 0 , 0 , n86 );
and_AQFP n87_( clk_8 , buf_N74_n87_3 , splitterfromn86 , 0 , 0 , n87 );
and_AQFP n88_( clk_3 , splittern83ton179n88 , buf_n87_n88_1 , 0 , 0 , n88 );
and_AQFP n89_( clk_7 , buf_N89_n89_2 , buf_splitterfromn78_n89_1 , 0 , 0 , n89 );
or_AQFP n90_( clk_4 , splitterN130ton120n91 , splitterN96ton273n91 , 0 , 0 , n90 );
and_AQFP n91_( clk_4 , splitterN130ton120n91 , splitterN96ton273n91 , 0 , 0 , n91 );
and_AQFP n92_( clk_5 , n90 , n91 , 0 , 1 , n92 );
and_AQFP n93_( clk_8 , splitterN91ton262n94 , splitterfromn92 , 0 , 0 , n93 );
or_AQFP n94_( clk_8 , splitterN91ton262n94 , splitterfromn92 , 0 , 0 , n94 );
and_AQFP n95_( clk_4 , buf_n93_n95_1 , buf_n94_n95_1 , 1 , 0 , n95 );
or_AQFP n96_( clk_6 , splitterN121ton182n97 , splitterfromN135 , 0 , 0 , n96 );
and_AQFP n97_( clk_6 , splitterN121ton182n97 , splitterfromN135 , 0 , 0 , n97 );
and_AQFP n98_( clk_7 , n96 , n97 , 0 , 1 , n98 );
and_AQFP n99_( clk_1 , splitterN126ton100n99 , splitterfromn98 , 0 , 1 , n99 );
and_AQFP n100_( clk_1 , splitterN126ton100n99 , splitterfromn98 , 1 , 0 , n100 );
or_AQFP n101_( clk_2 , n99 , n100 , 0 , 0 , n101 );
and_AQFP n102_( clk_6 , splitterN101ton102n316 , splitterN106ton102n289 , 0 , 1 , n102 );
and_AQFP n103_( clk_6 , splitterN101ton102n316 , splitterN106ton102n289 , 1 , 0 , n103 );
or_AQFP n104_( clk_7 , n102 , n103 , 0 , 0 , n104 );
or_AQFP n105_( clk_6 , splitterN111ton105n237 , splitterN116ton105n255 , 0 , 0 , n105 );
and_AQFP n106_( clk_6 , splitterN111ton105n237 , splitterN116ton105n255 , 0 , 0 , n106 );
and_AQFP n107_( clk_7 , n105 , n106 , 0 , 1 , n107 );
or_AQFP n108_( clk_2 , splitterfromn104 , splitterfromn107 , 0 , 0 , n108 );
and_AQFP n109_( clk_3 , buf_splitterfromn104_n109_1 , splitterfromn107 , 0 , 0 , n109 );
and_AQFP n110_( clk_4 , n108 , n109 , 0 , 1 , n110 );
or_AQFP n111_( clk_6 , splitterfromn101 , splitterfromn110 , 0 , 0 , n111 );
and_AQFP n112_( clk_6 , splitterfromn101 , splitterfromn110 , 0 , 0 , n112 );
and_AQFP n113_( clk_8 , n111 , n112 , 0 , 1 , n113 );
and_AQFP n114_( clk_1 , buf_splitterfromn95_n114_12 , buf_splitterfromn113_n114_13 , 1 , 0 , n114 );
and_AQFP n115_( clk_8 , buf_splitterfromn95_n115_8 , buf_splitterfromn113_n115_5 , 0 , 1 , n115 );
or_AQFP n116_( clk_2 , n114 , buf_n115_n116_4 , 0 , 0 , n116 );
or_AQFP n117_( clk_6 , splitterN159ton117n330 , splitterN177ton117n315 , 0 , 0 , n117 );
and_AQFP n118_( clk_6 , splitterN159ton117n330 , splitterN177ton117n315 , 0 , 0 , n118 );
and_AQFP n119_( clk_8 , n117 , n118 , 0 , 1 , n119 );
and_AQFP n120_( clk_4 , buf_splitterN130ton120n91_n120_4 , splitterfromn119 , 0 , 1 , n120 );
and_AQFP n121_( clk_4 , buf_splitterN130ton120n91_n121_4 , splitterfromn119 , 1 , 0 , n121 );
or_AQFP n122_( clk_6 , n120 , n121 , 0 , 0 , n122 );
or_AQFP n123_( clk_1 , buf_splitterN189ton123n236_n123_1 , splitterN195ton123n253 , 0 , 0 , n123 );
and_AQFP n124_( clk_2 , buf_splitterN189ton123n236_n124_2 , buf_splitterN195ton123n253_n124_1 , 0 , 0 , n124 );
and_AQFP n125_( clk_3 , n123 , n124 , 0 , 1 , n125 );
and_AQFP n126_( clk_5 , splitterfromN207 , splitterfromn125 , 0 , 1 , n126 );
and_AQFP n127_( clk_5 , splitterfromN207 , splitterfromn125 , 1 , 0 , n127 );
or_AQFP n128_( clk_6 , n126 , n127 , 0 , 0 , n128 );
and_AQFP n129_( clk_7 , splitterN165ton129n346 , splitterN201ton129n180 , 1 , 0 , n129 );
and_AQFP n130_( clk_7 , splitterN165ton129n346 , splitterN201ton129n180 , 0 , 1 , n130 );
or_AQFP n131_( clk_1 , n129 , n130 , 0 , 0 , n131 );
and_AQFP n132_( clk_1 , splitterN171ton132n361 , splitterN183ton132n221 , 0 , 1 , n132 );
and_AQFP n133_( clk_1 , splitterN171ton132n361 , splitterN183ton132n221 , 1 , 0 , n133 );
or_AQFP n134_( clk_2 , n132 , n133 , 0 , 0 , n134 );
and_AQFP n135_( clk_5 , splitterfromn131 , splitterfromn134 , 0 , 1 , n135 );
and_AQFP n136_( clk_5 , buf_splitterfromn131_n136_1 , buf_splitterfromn134_n136_1 , 1 , 0 , n136 );
or_AQFP n137_( clk_7 , n135 , n136 , 0 , 0 , n137 );
and_AQFP n138_( clk_2 , splitterfromn128 , splitterfromn137 , 1 , 0 , n138 );
and_AQFP n139_( clk_2 , splitterfromn128 , splitterfromn137 , 0 , 1 , n139 );
or_AQFP n140_( clk_4 , n138 , n139 , 0 , 0 , n140 );
and_AQFP n141_( clk_2 , buf_splitterfromn122_n141_1 , splitterfromn140 , 0 , 1 , n141 );
and_AQFP n142_( clk_3 , buf_splitterfromn122_n142_3 , splitterfromn140 , 1 , 0 , n142 );
or_AQFP n143_( clk_4 , n141 , n142 , 0 , 0 , n143 );
and_AQFP n144_( clk_3 , N156 , splitterN59ton144n86 , 0 , 0 , n144 );
and_AQFP n145_( clk_7 , splittern81toN447n156 , buf_splitterfromn144_n145_1 , 0 , 1 , n145 );
and_AQFP n146_( clk_1 , buf_splitterN17ton146n68_n146_3 , splitterfromn145 , 0 , 0 , n146 );
and_AQFP n147_( clk_2 , buf_splitterN1ton147n70_n147_4 , n146 , 0 , 1 , n147 );
and_AQFP n148_( clk_4 , buf_splitterfromN153_n148_2 , splittern147ton148n208 , 0 , 1 , n148 );
and_AQFP n149_( clk_6 , splitterN80ton149n76 , splitterfromn61 , 0 , 0 , n149 );
and_AQFP n150_( clk_7 , splittern81toN447n156 , n149 , 0 , 0 , n150 );
and_AQFP n151_( clk_1 , buf_splitterN55ton151n82_n151_1 , splitterfromn150 , 0 , 0 , n151 );
and_AQFP n152_( clk_2 , buf_splitterN268ton152n331_n152_2 , n151 , 1 , 0 , n152 );
and_AQFP n153_( clk_4 , splitterN17ton146n68 , splitterN42ton153n77 , 0 , 1 , n153 );
and_AQFP n154_( clk_4 , splitterN17ton146n68 , splitterN42ton153n77 , 1 , 0 , n154 );
or_AQFP n155_( clk_7 , buf_n153_n155_1 , buf_n154_n155_1 , 0 , 0 , n155 );
and_AQFP n156_( clk_7 , splittern81toN447n156 , buf_splitterfromn144_n156_1 , 0 , 0 , n156 );
and_AQFP n157_( clk_8 , n155 , n156 , 0 , 0 , n157 );
and_AQFP n158_( clk_7 , buf_splitterN42ton153n77_n158_1 , splitterfromn73 , 0 , 0 , n158 );
and_AQFP n159_( clk_5 , splitterN17ton159n68 , splitterN51ton159n81 , 0 , 0 , n159 );
and_AQFP n160_( clk_7 , splittern67ton160n83 , n159 , 0 , 0 , n160 );
and_AQFP n161_( clk_8 , n158 , n160 , 1 , 0 , n161 );
or_AQFP n162_( clk_1 , n157 , n161 , 0 , 0 , n162 );
and_AQFP n163_( clk_3 , buf_splitterN126ton100n99_n163_1 , splittern162ton163n289 , 0 , 0 , n163 );
or_AQFP n164_( clk_4 , splittern152ton164n210 , n163 , 0 , 0 , n164 );
or_AQFP n165_( clk_5 , n148 , n164 , 0 , 0 , n165 );
or_AQFP n166_( clk_7 , buf_splitterN201ton129n180_n166_4 , splittern165ton166n175 , 0 , 0 , n166 );
and_AQFP n167_( clk_7 , buf_splitterN201ton167n180_n167_3 , splittern165ton166n175 , 0 , 0 , n167 );
and_AQFP n168_( clk_1 , splitterfromn166 , splittern167ton168n201 , 0 , 1 , n168 );
and_AQFP n169_( clk_3 , buf_splitterN261ton169n201_n169_3 , splittern168ton169n173 , 0 , 0 , n169 );
or_AQFP n170_( clk_3 , buf_splitterN261ton169n201_n170_3 , splittern168ton169n173 , 0 , 0 , n170 );
and_AQFP n171_( clk_4 , buf_splitterN219ton171n355_n171_3 , n170 , 0 , 0 , n171 );
and_AQFP n172_( clk_5 , n169 , n171 , 1 , 0 , n172 );
and_AQFP n173_( clk_3 , buf_splitterN228ton173n357_n173_3 , splittern168ton169n173 , 0 , 0 , n173 );
and_AQFP n174_( clk_1 , buf_splitterN237ton174n358_n174_5 , splittern167ton168n201 , 0 , 0 , n174 );
and_AQFP n175_( clk_7 , buf_splitterN246ton175n359_n175_1 , splittern165ton166n175 , 0 , 0 , n175 );
and_AQFP n176_( clk_6 , splitterN42ton176n77 , buf_N72_n176_2 , 0 , 0 , n176 );
and_AQFP n177_( clk_7 , buf_N73_n177_2 , n176 , 0 , 0 , n177 );
and_AQFP n178_( clk_8 , splitterfromn86 , n177 , 0 , 0 , n178 );
and_AQFP n179_( clk_2 , splittern83ton179n88 , n178 , 0 , 0 , n179 );
and_AQFP n180_( clk_4 , splitterN201ton167n180 , splittern179ton180n361 , 0 , 0 , n180 );
and_AQFP n181_( clk_7 , splitterN255ton181n254 , buf_N267_n181_2 , 0 , 0 , n181 );
and_AQFP n182_( clk_7 , splitterN121ton182n97 , buf_splitterN210ton182n360_n182_1 , 0 , 0 , n182 );
or_AQFP n183_( clk_3 , buf_n181_n183_2 , buf_n182_n183_1 , 0 , 0 , n183 );
or_AQFP n184_( clk_6 , n180 , buf_n183_n184_1 , 0 , 0 , n184 );
or_AQFP n185_( clk_1 , n175 , buf_n184_n185_1 , 0 , 0 , n185 );
or_AQFP n186_( clk_2 , n174 , n185 , 0 , 0 , n186 );
or_AQFP n187_( clk_4 , n173 , n186 , 0 , 0 , n187 );
or_AQFP n188_( clk_7 , n172 , buf_n187_n188_1 , 0 , 0 , n188 );
and_AQFP n189_( clk_4 , buf_splitterfromN146_n189_2 , splittern147ton148n208 , 0 , 1 , n189 );
and_AQFP n190_( clk_3 , buf_splitterN116ton105n255_n190_2 , splittern162ton163n289 , 0 , 0 , n190 );
or_AQFP n191_( clk_4 , splittern152ton164n210 , n190 , 0 , 0 , n191 );
or_AQFP n192_( clk_5 , n189 , n191 , 0 , 0 , n192 );
and_AQFP n193_( clk_7 , buf_splitterN189ton123n236_n193_4 , splittern192ton193n235 , 0 , 0 , n193 );
or_AQFP n194_( clk_7 , splitterN189ton194n236 , splittern192ton193n235 , 0 , 0 , n194 );
and_AQFP n195_( clk_4 , splitterfromN149 , splittern147ton148n208 , 0 , 1 , n195 );
and_AQFP n196_( clk_4 , buf_splitterN121ton182n97_n196_3 , splittern162ton196n207 , 0 , 0 , n196 );
or_AQFP n197_( clk_5 , splittern152ton164n210 , n196 , 0 , 0 , n197 );
or_AQFP n198_( clk_6 , n195 , n197 , 0 , 0 , n198 );
and_AQFP n199_( clk_8 , buf_splitterN195ton123n253_n199_3 , splittern198ton199n252 , 0 , 0 , n199 );
or_AQFP n200_( clk_8 , buf_splitterN195ton200n253_n200_3 , splittern198ton199n252 , 0 , 0 , n200 );
or_AQFP n201_( clk_1 , buf_splitterN261ton169n201_n201_2 , splittern167ton168n201 , 0 , 0 , n201 );
and_AQFP n202_( clk_2 , splitterfromn166 , n201 , 0 , 0 , n202 );
and_AQFP n203_( clk_4 , buf_splitterfromn200_n203_1 , splittern202ton203n247 , 0 , 0 , n203 );
or_AQFP n204_( clk_5 , buf_splittern199ton204n251_n204_1 , n203 , 0 , 0 , n204 );
and_AQFP n205_( clk_7 , buf_splitterfromn194_n205_3 , splittern204ton205n230 , 0 , 0 , n205 );
or_AQFP n206_( clk_8 , buf_splittern193ton206n234_n206_4 , n205 , 0 , 0 , n206 );
and_AQFP n207_( clk_4 , buf_splitterN111ton105n237_n207_3 , splittern162ton196n207 , 0 , 0 , n207 );
and_AQFP n208_( clk_4 , splitterfromN143 , splittern147ton148n208 , 0 , 1 , n208 );
or_AQFP n209_( clk_5 , n207 , n208 , 0 , 0 , n209 );
or_AQFP n210_( clk_6 , buf_splittern152ton164n210_n210_2 , n209 , 0 , 0 , n210 );
and_AQFP n211_( clk_8 , buf_splitterN183ton132n221_n211_3 , splittern210ton211n220 , 0 , 0 , n211 );
or_AQFP n212_( clk_8 , buf_splitterN183ton212n221_n212_3 , splittern210ton211n220 , 0 , 0 , n212 );
and_AQFP n213_( clk_2 , splittern211ton213n298 , splitterfromn212 , 1 , 0 , n213 );
or_AQFP n214_( clk_2 , splittern206ton214n297 , buf_splittern213ton214n218_n214_3 , 0 , 0 , n214 );
and_AQFP n215_( clk_2 , splittern206ton214n297 , buf_splittern213ton214n218_n215_3 , 0 , 0 , n215 );
and_AQFP n216_( clk_3 , n214 , n215 , 0 , 1 , n216 );
and_AQFP n217_( clk_5 , buf_splitterN219ton171n355_n217_7 , n216 , 0 , 0 , n217 );
and_AQFP n218_( clk_4 , buf_splitterN228ton173n357_n218_2 , splittern213ton214n218 , 0 , 0 , n218 );
and_AQFP n219_( clk_3 , buf_splitterN237ton174n358_n219_6 , splittern211ton213n298 , 0 , 0 , n219 );
and_AQFP n220_( clk_8 , buf_splitterN246ton175n359_n220_1 , splittern210ton211n220 , 0 , 0 , n220 );
and_AQFP n221_( clk_5 , splitterN183ton212n221 , splittern179ton180n361 , 0 , 0 , n221 );
and_AQFP n222_( clk_7 , splitterN106ton102n289 , splitterN210ton182n360 , 0 , 0 , n222 );
or_AQFP n223_( clk_6 , n221 , buf_n222_n223_3 , 0 , 0 , n223 );
or_AQFP n224_( clk_2 , n220 , buf_n223_n224_3 , 0 , 0 , n224 );
or_AQFP n225_( clk_5 , n219 , buf_n224_n225_1 , 0 , 0 , n225 );
or_AQFP n226_( clk_3 , buf_n218_n226_3 , buf_n225_n226_2 , 0 , 0 , n226 );
or_AQFP n227_( clk_6 , buf_n217_n227_5 , buf_n226_n227_6 , 0 , 0 , n227 );
and_AQFP n228_( clk_1 , splittern193ton206n234 , splitterfromn194 , 1 , 0 , n228 );
or_AQFP n229_( clk_7 , splittern204ton205n230 , buf_splittern228ton229n233_n229_2 , 0 , 0 , n229 );
and_AQFP n230_( clk_7 , splittern204ton205n230 , buf_splittern228ton229n233_n230_2 , 0 , 0 , n230 );
and_AQFP n231_( clk_8 , n229 , n230 , 0 , 1 , n231 );
and_AQFP n232_( clk_1 , buf_splitterN219ton232n308_n232_1 , n231 , 0 , 0 , n232 );
and_AQFP n233_( clk_3 , splitterN228ton233n250 , splittern228ton229n233 , 0 , 0 , n233 );
and_AQFP n234_( clk_1 , splitterN237ton234n251 , splittern193ton206n234 , 0 , 0 , n234 );
and_AQFP n235_( clk_7 , splitterN246ton235n252 , splittern192ton193n235 , 0 , 0 , n235 );
and_AQFP n236_( clk_6 , splitterN189ton194n236 , splittern179ton236n253 , 0 , 0 , n236 );
and_AQFP n237_( clk_7 , splitterN111ton105n237 , splitterN210ton237n255 , 0 , 0 , n237 );
and_AQFP n238_( clk_6 , splitterN255ton181n254 , buf_N259_n238_2 , 0 , 0 , n238 );
or_AQFP n239_( clk_2 , buf_n237_n239_1 , buf_n238_n239_3 , 0 , 0 , n239 );
or_AQFP n240_( clk_7 , n236 , buf_n239_n240_4 , 0 , 0 , n240 );
or_AQFP n241_( clk_1 , n235 , n240 , 0 , 0 , n241 );
or_AQFP n242_( clk_2 , n234 , n241 , 0 , 0 , n242 );
or_AQFP n243_( clk_4 , n233 , n242 , 0 , 0 , n243 );
or_AQFP n244_( clk_2 , n232 , buf_n243_n244_3 , 0 , 0 , n244 );
and_AQFP n245_( clk_2 , splittern199ton204n251 , splitterfromn200 , 1 , 0 , n245 );
or_AQFP n246_( clk_4 , splittern202ton203n247 , splittern245ton246n250 , 0 , 0 , n246 );
and_AQFP n247_( clk_4 , splittern202ton203n247 , splittern245ton246n250 , 0 , 0 , n247 );
and_AQFP n248_( clk_5 , n246 , n247 , 0 , 1 , n248 );
and_AQFP n249_( clk_6 , splitterN219ton232n308 , n248 , 0 , 0 , n249 );
and_AQFP n250_( clk_4 , splitterN228ton233n250 , splittern245ton246n250 , 0 , 0 , n250 );
and_AQFP n251_( clk_2 , splitterN237ton234n251 , splittern199ton204n251 , 0 , 0 , n251 );
and_AQFP n252_( clk_8 , splitterN246ton235n252 , splittern198ton199n252 , 0 , 0 , n252 );
and_AQFP n253_( clk_7 , buf_splitterN195ton200n253_n253_1 , splittern179ton236n253 , 0 , 0 , n253 );
and_AQFP n254_( clk_7 , splitterN255ton181n254 , buf_N260_n254_2 , 0 , 0 , n254 );
and_AQFP n255_( clk_8 , buf_splitterN116ton105n255_n255_1 , splitterN210ton237n255 , 0 , 0 , n255 );
or_AQFP n256_( clk_1 , n254 , n255 , 0 , 0 , n256 );
or_AQFP n257_( clk_1 , n253 , buf_n256_n257_5 , 0 , 0 , n257 );
or_AQFP n258_( clk_2 , n252 , n257 , 0 , 0 , n258 );
or_AQFP n259_( clk_3 , n251 , n258 , 0 , 0 , n259 );
or_AQFP n260_( clk_5 , n250 , buf_n259_n260_1 , 0 , 0 , n260 );
or_AQFP n261_( clk_7 , n249 , n260 , 0 , 0 , n261 );
and_AQFP n262_( clk_4 , buf_splitterN91ton262n94_n262_2 , splittern162ton262n289 , 0 , 0 , n262 );
and_AQFP n263_( clk_1 , buf_splitterN55ton151n82_n263_2 , splitterfromn145 , 0 , 0 , n263 );
and_AQFP n264_( clk_3 , splitterfromN143 , splittern263ton264n290 , 0 , 0 , n264 );
and_AQFP n265_( clk_5 , splitterN17ton159n68 , splitterN268ton152n331 , 0 , 1 , n265 );
and_AQFP n266_( clk_1 , splitterfromn150 , buf_n265_n266_1 , 0 , 0 , n266 );
and_AQFP n267_( clk_2 , buf_splitterN138ton267n291_n267_1 , buf_splitterfromN8_n267_4 , 0 , 0 , n267 );
or_AQFP n268_( clk_3 , splittern266ton268n292 , n267 , 0 , 0 , n268 );
or_AQFP n269_( clk_4 , n264 , n268 , 0 , 0 , n269 );
or_AQFP n270_( clk_5 , n262 , n269 , 0 , 0 , n270 );
and_AQFP n271_( clk_7 , buf_splitterN159ton117n330_n271_5 , splittern270ton271n329 , 0 , 0 , n271 );
or_AQFP n272_( clk_7 , splitterN159ton272n330 , splittern270ton271n329 , 0 , 0 , n272 );
and_AQFP n273_( clk_4 , buf_splitterN96ton273n91_n273_5 , splittern162ton262n289 , 0 , 0 , n273 );
and_AQFP n274_( clk_3 , buf_splitterfromN146_n274_1 , splittern263ton264n290 , 0 , 0 , n274 );
and_AQFP n275_( clk_1 , splitterN138ton267n291 , buf_splitterN51ton159n81_n275_2 , 0 , 0 , n275 );
or_AQFP n276_( clk_3 , splittern266ton268n292 , n275 , 0 , 0 , n276 );
or_AQFP n277_( clk_4 , n274 , n276 , 0 , 0 , n277 );
or_AQFP n278_( clk_5 , n273 , n277 , 0 , 0 , n278 );
and_AQFP n279_( clk_7 , buf_splitterN165ton129n346_n279_5 , splittern278ton279n344 , 0 , 0 , n279 );
or_AQFP n280_( clk_8 , buf_splitterN165ton280n346_n280_1 , splittern278ton279n344 , 0 , 0 , n280 );
and_AQFP n281_( clk_4 , buf_splitterN101ton102n316_n281_3 , splittern162ton262n289 , 0 , 0 , n281 );
and_AQFP n282_( clk_3 , splitterfromN149 , splittern263ton264n290 , 0 , 0 , n282 );
and_AQFP n283_( clk_2 , buf_splitterN138ton267n291_n283_1 , buf_splitterN17ton159n68_n283_3 , 0 , 0 , n283 );
or_AQFP n284_( clk_3 , splittern266ton268n292 , n283 , 0 , 0 , n284 );
or_AQFP n285_( clk_4 , n282 , n284 , 0 , 0 , n285 );
or_AQFP n286_( clk_5 , n281 , n285 , 0 , 0 , n286 );
and_AQFP n287_( clk_7 , buf_splitterN171ton132n361_n287_3 , splittern286ton287n359 , 0 , 0 , n287 );
or_AQFP n288_( clk_7 , buf_splitterN171ton288n361_n288_1 , splittern286ton287n359 , 0 , 0 , n288 );
and_AQFP n289_( clk_4 , buf_splitterN106ton102n289_n289_3 , splittern162ton262n289 , 0 , 0 , n289 );
and_AQFP n290_( clk_3 , buf_splitterfromN153_n290_2 , splittern263ton264n290 , 0 , 0 , n290 );
and_AQFP n291_( clk_1 , splitterN138ton267n291 , buf_N152_n291_3 , 0 , 0 , n291 );
or_AQFP n292_( clk_3 , splittern266ton268n292 , n291 , 0 , 0 , n292 );
or_AQFP n293_( clk_4 , n290 , n292 , 0 , 0 , n293 );
or_AQFP n294_( clk_5 , n289 , n293 , 0 , 0 , n294 );
and_AQFP n295_( clk_7 , buf_splitterN177ton117n315_n295_4 , splittern294ton295n314 , 0 , 0 , n295 );
or_AQFP n296_( clk_8 , buf_splitterN177ton296n315_n296_2 , splittern294ton295n314 , 0 , 0 , n296 );
and_AQFP n297_( clk_2 , splittern206ton214n297 , buf_splitterfromn212_n297_6 , 0 , 0 , n297 );
or_AQFP n298_( clk_3 , buf_splittern211ton213n298_n298_4 , n297 , 0 , 0 , n298 );
and_AQFP n299_( clk_5 , buf_splitterfromn296_n299_5 , splittern298ton299n312 , 0 , 0 , n299 );
or_AQFP n300_( clk_6 , buf_splittern295ton300n313_n300_6 , n299 , 0 , 0 , n300 );
and_AQFP n301_( clk_8 , buf_splitterfromn288_n301_8 , splittern300ton301n354 , 0 , 0 , n301 );
or_AQFP n302_( clk_1 , buf_splittern287ton302n358_n302_9 , n301 , 0 , 0 , n302 );
and_AQFP n303_( clk_3 , buf_splitterfromn280_n303_5 , splittern302ton303n339 , 0 , 0 , n303 );
or_AQFP n304_( clk_4 , buf_splittern279ton304n343_n304_9 , n303 , 0 , 0 , n304 );
and_AQFP n305_( clk_6 , buf_splitterfromn272_n305_10 , splittern304ton305n324 , 0 , 0 , n305 );
or_AQFP n306_( clk_8 , buf_splittern271ton306n328_n306_12 , n305 , 0 , 0 , n306 );
and_AQFP n307_( clk_4 , buf_splittern295ton300n313_n307_1 , splitterfromn296 , 1 , 0 , n307 );
and_AQFP n308_( clk_5 , buf_splitterN219ton232n308_n308_4 , splittern298ton299n312 , 0 , 1 , n308 );
or_AQFP n309_( clk_7 , buf_splitterN228ton309n357_n309_5 , n308 , 0 , 0 , n309 );
and_AQFP n310_( clk_8 , buf_splitterfromn307_n310_3 , n309 , 0 , 0 , n310 );
and_AQFP n311_( clk_6 , splitterN219ton311n355 , buf_splitterfromn307_n311_2 , 0 , 1 , n311 );
and_AQFP n312_( clk_7 , buf_splittern298ton299n312_n312_1 , n311 , 0 , 0 , n312 );
and_AQFP n313_( clk_2 , buf_splitterN237ton313n358_n313_1 , splittern295ton300n313 , 0 , 0 , n313 );
and_AQFP n314_( clk_7 , splitterN246ton314n359 , splittern294ton295n314 , 0 , 0 , n314 );
and_AQFP n315_( clk_6 , splitterN177ton296n315 , splittern179ton315n361 , 0 , 0 , n315 );
and_AQFP n316_( clk_8 , buf_splitterN101ton102n316_n316_1 , splitterN210ton316n360 , 0 , 0 , n316 );
or_AQFP n317_( clk_7 , n315 , buf_n316_n317_3 , 0 , 0 , n317 );
or_AQFP n318_( clk_8 , n314 , n317 , 0 , 0 , n318 );
or_AQFP n319_( clk_3 , n313 , buf_n318_n319_1 , 0 , 0 , n319 );
or_AQFP n320_( clk_8 , n312 , buf_n319_n320_8 , 0 , 0 , n320 );
or_AQFP n321_( clk_2 , n310 , n320 , 0 , 0 , n321 );
and_AQFP n322_( clk_2 , splittern271ton306n328 , splitterfromn272 , 1 , 0 , n322 );
or_AQFP n323_( clk_6 , splittern304ton305n324 , buf_splittern322ton323n327_n323_9 , 0 , 0 , n323 );
and_AQFP n324_( clk_7 , splittern304ton305n324 , buf_splittern322ton323n327_n324_10 , 0 , 0 , n324 );
and_AQFP n325_( clk_8 , buf_splitterN219ton311n355_n325_6 , n324 , 0 , 1 , n325 );
and_AQFP n326_( clk_1 , buf_n323_n326_1 , n325 , 0 , 0 , n326 );
and_AQFP n327_( clk_5 , splitterN228ton309n357 , splittern322ton323n327 , 0 , 0 , n327 );
and_AQFP n328_( clk_1 , buf_splitterN237ton313n358_n328_1 , splittern271ton306n328 , 0 , 0 , n328 );
and_AQFP n329_( clk_7 , splitterN246ton314n359 , splittern270ton271n329 , 0 , 0 , n329 );
and_AQFP n330_( clk_6 , splitterN159ton272n330 , splittern179ton315n361 , 0 , 0 , n330 );
and_AQFP n331_( clk_8 , splitterN210ton316n360 , buf_splitterN268ton152n331_n331_1 , 0 , 0 , n331 );
or_AQFP n332_( clk_7 , n330 , buf_n331_n332_3 , 0 , 0 , n332 );
or_AQFP n333_( clk_8 , n329 , n332 , 0 , 0 , n333 );
or_AQFP n334_( clk_2 , n328 , n333 , 0 , 0 , n334 );
or_AQFP n335_( clk_1 , buf_n327_n335_1 , buf_n334_n335_4 , 0 , 0 , n335 );
or_AQFP n336_( clk_3 , n326 , buf_n335_n336_12 , 0 , 0 , n336 );
and_AQFP n337_( clk_8 , buf_splittern279ton304n343_n337_3 , splitterfromn280 , 1 , 0 , n337 );
and_AQFP n338_( clk_4 , splittern302ton303n339 , buf_splittern337ton338n342_n338_3 , 0 , 0 , n338 );
or_AQFP n339_( clk_4 , splittern302ton303n339 , buf_splittern337ton338n342_n339_5 , 0 , 0 , n339 );
and_AQFP n340_( clk_5 , buf_splitterN219ton311n355_n340_4 , n339 , 0 , 0 , n340 );
and_AQFP n341_( clk_6 , n338 , n340 , 1 , 0 , n341 );
and_AQFP n342_( clk_8 , buf_splitterN228ton309n357_n342_11 , splittern337ton338n342 , 0 , 0 , n342 );
and_AQFP n343_( clk_1 , buf_splitterN237ton313n358_n343_1 , splittern279ton304n343 , 0 , 0 , n343 );
and_AQFP n344_( clk_7 , splitterN246ton314n359 , splittern278ton279n344 , 0 , 0 , n344 );
and_AQFP n345_( clk_1 , splitterN210ton316n360 , buf_splitterN91ton262n94_n345_2 , 0 , 0 , n345 );
and_AQFP n346_( clk_6 , splitterN165ton280n346 , splittern179ton315n361 , 0 , 0 , n346 );
or_AQFP n347_( clk_7 , buf_n345_n347_3 , n346 , 0 , 0 , n347 );
or_AQFP n348_( clk_8 , n344 , n347 , 0 , 0 , n348 );
or_AQFP n349_( clk_2 , n343 , n348 , 0 , 0 , n349 );
or_AQFP n350_( clk_1 , n342 , buf_n349_n350_12 , 0 , 0 , n350 );
or_AQFP n351_( clk_8 , n341 , buf_n350_n351_6 , 0 , 0 , n351 );
and_AQFP n352_( clk_2 , splittern287ton302n358 , splitterfromn288 , 1 , 0 , n352 );
and_AQFP n353_( clk_8 , splittern300ton301n354 , buf_splittern352ton353n357_n353_7 , 0 , 0 , n353 );
or_AQFP n354_( clk_8 , splittern300ton301n354 , buf_splittern352ton353n357_n354_6 , 0 , 0 , n354 );
and_AQFP n355_( clk_1 , buf_splitterN219ton311n355_n355_2 , n354 , 0 , 0 , n355 );
and_AQFP n356_( clk_2 , n353 , n355 , 1 , 0 , n356 );
and_AQFP n357_( clk_6 , buf_splitterN228ton309n357_n357_1 , splittern352ton353n357 , 0 , 0 , n357 );
and_AQFP n358_( clk_1 , buf_splitterN237ton313n358_n358_2 , splittern287ton302n358 , 0 , 0 , n358 );
and_AQFP n359_( clk_7 , splitterN246ton314n359 , splittern286ton287n359 , 0 , 0 , n359 );
and_AQFP n360_( clk_1 , splitterN210ton316n360 , buf_splitterN96ton273n91_n360_2 , 0 , 0 , n360 );
and_AQFP n361_( clk_5 , splitterN171ton288n361 , splittern179ton315n361 , 0 , 0 , n361 );
or_AQFP n362_( clk_6 , buf_n360_n362_4 , n361 , 0 , 0 , n362 );
or_AQFP n363_( clk_8 , n359 , buf_n362_n363_1 , 0 , 0 , n363 );
or_AQFP n364_( clk_2 , n358 , n363 , 0 , 0 , n364 );
or_AQFP n365_( clk_8 , n357 , buf_n364_n365_5 , 0 , 0 , n365 );
or_AQFP n366_( clk_1 , buf_n356_n366_3 , buf_n365_n366_11 , 0 , 0 , n366 );
PO_AQFP N388_( clk_5 , buf_n62_N388_18 , 0 , N388 );
PO_AQFP N389_( clk_5 , buf_n64_N389_18 , 0 , N389 );
PO_AQFP N390_( clk_5 , buf_splittern65toN390n80_N390_1 , 0 , N390 );
PO_AQFP N391_( clk_5 , buf_n66_N391_21 , 0 , N391 );
PO_AQFP N418_( clk_5 , buf_n69_N418_7 , 0 , N418 );
PO_AQFP N419_( clk_5 , buf_n72_N419_1 , 1 , N419 );
PO_AQFP N420_( clk_5 , buf_n74_N420_18 , 1 , N420 );
PO_AQFP N421_( clk_5 , buf_n76_N421_9 , 1 , N421 );
PO_AQFP N422_( clk_5 , buf_n77_N422_24 , 1 , N422 );
PO_AQFP N423_( clk_5 , buf_n79_N423_21 , 0 , N423 );
PO_AQFP N446_( clk_5 , buf_n80_N446_1 , 1 , N446 );
PO_AQFP N447_( clk_5 , buf_splittern81toN447n156_N447_19 , 0 , N447 );
PO_AQFP N448_( clk_5 , buf_n85_N448_3 , 0 , N448 );
PO_AQFP N449_( clk_5 , buf_n88_N449_17 , 0 , N449 );
PO_AQFP N450_( clk_5 , buf_n89_N450_36 , 0 , N450 );
PO_AQFP N767_( clk_5 , buf_n116_N767_1 , 0 , N767 );
PO_AQFP N768_( clk_5 , buf_n143_N768_10 , 0 , N768 );
PO_AQFP N850_( clk_5 , buf_n188_N850_12 , 0 , N850 );
PO_AQFP N863_( clk_5 , buf_n227_N863_6 , 0 , N863 );
PO_AQFP N864_( clk_5 , buf_n244_N864_15 , 0 , N864 );
PO_AQFP N865_( clk_5 , buf_n261_N865_11 , 0 , N865 );
PO_AQFP N866_( clk_5 , buf_n306_N866_2 , 0 , N866 );
PO_AQFP N874_( clk_5 , buf_n321_N874_7 , 0 , N874 );
PO_AQFP N878_( clk_5 , n336 , 0 , N878 );
PO_AQFP N879_( clk_5 , buf_n351_N879_2 , 0 , N879 );
PO_AQFP N880_( clk_5 , buf_n366_N880_1 , 0 , N880 );
buf_AQFP buf_N101_splitterN101ton102n316_1_( clk_3 , N101 , 0 , buf_N101_splitterN101ton102n316_1 );
buf_AQFP buf_N106_splitterN106ton102n289_1_( clk_3 , N106 , 0 , buf_N106_splitterN106ton102n289_1 );
buf_AQFP buf_N111_splitterN111ton105n237_1_( clk_3 , N111 , 0 , buf_N111_splitterN111ton105n237_1 );
buf_AQFP buf_N116_splitterN116ton105n255_1_( clk_3 , N116 , 0 , buf_N116_splitterN116ton105n255_1 );
buf_AQFP buf_N121_splitterN121ton182n97_1_( clk_3 , N121 , 0 , buf_N121_splitterN121ton182n97_1 );
buf_AQFP buf_N121_splitterN121ton182n97_2_( clk_4 , buf_N121_splitterN121ton182n97_1 , 0 , buf_N121_splitterN121ton182n97_2 );
buf_AQFP buf_N126_splitterN126ton100n99_1_( clk_3 , N126 , 0 , buf_N126_splitterN126ton100n99_1 );
buf_AQFP buf_N126_splitterN126ton100n99_2_( clk_5 , buf_N126_splitterN126ton100n99_1 , 0 , buf_N126_splitterN126ton100n99_2 );
buf_AQFP buf_N13_splitterfromN13_1_( clk_3 , N13 , 0 , buf_N13_splitterfromN13_1 );
buf_AQFP buf_N135_splitterfromN135_1_( clk_3 , N135 , 0 , buf_N135_splitterfromN135_1 );
buf_AQFP buf_N138_splitterN138ton267n291_1_( clk_3 , N138 , 0 , buf_N138_splitterN138ton267n291_1 );
buf_AQFP buf_N138_splitterN138ton267n291_2_( clk_5 , buf_N138_splitterN138ton267n291_1 , 0 , buf_N138_splitterN138ton267n291_2 );
buf_AQFP buf_N143_splitterfromN143_1_( clk_3 , N143 , 0 , buf_N143_splitterfromN143_1 );
buf_AQFP buf_N143_splitterfromN143_2_( clk_4 , buf_N143_splitterfromN143_1 , 0 , buf_N143_splitterfromN143_2 );
buf_AQFP buf_N143_splitterfromN143_3_( clk_5 , buf_N143_splitterfromN143_2 , 0 , buf_N143_splitterfromN143_3 );
buf_AQFP buf_N143_splitterfromN143_4_( clk_7 , buf_N143_splitterfromN143_3 , 0 , buf_N143_splitterfromN143_4 );
buf_AQFP buf_N143_splitterfromN143_5_( clk_8 , buf_N143_splitterfromN143_4 , 0 , buf_N143_splitterfromN143_5 );
buf_AQFP buf_N146_splitterfromN146_1_( clk_3 , N146 , 0 , buf_N146_splitterfromN146_1 );
buf_AQFP buf_N146_splitterfromN146_2_( clk_5 , buf_N146_splitterfromN146_1 , 0 , buf_N146_splitterfromN146_2 );
buf_AQFP buf_N149_splitterfromN149_1_( clk_3 , N149 , 0 , buf_N149_splitterfromN149_1 );
buf_AQFP buf_N149_splitterfromN149_2_( clk_5 , buf_N149_splitterfromN149_1 , 0 , buf_N149_splitterfromN149_2 );
buf_AQFP buf_N149_splitterfromN149_3_( clk_7 , buf_N149_splitterfromN149_2 , 0 , buf_N149_splitterfromN149_3 );
buf_AQFP buf_N149_splitterfromN149_4_( clk_1 , buf_N149_splitterfromN149_3 , 0 , buf_N149_splitterfromN149_4 );
buf_AQFP buf_N152_n291_1_( clk_3 , N152 , 0 , buf_N152_n291_1 );
buf_AQFP buf_N152_n291_2_( clk_5 , buf_N152_n291_1 , 0 , buf_N152_n291_2 );
buf_AQFP buf_N152_n291_3_( clk_7 , buf_N152_n291_2 , 0 , buf_N152_n291_3 );
buf_AQFP buf_N153_splitterfromN153_1_( clk_3 , N153 , 0 , buf_N153_splitterfromN153_1 );
buf_AQFP buf_N153_splitterfromN153_2_( clk_5 , buf_N153_splitterfromN153_1 , 0 , buf_N153_splitterfromN153_2 );
buf_AQFP buf_N159_splitterN159ton117n330_1_( clk_3 , N159 , 0 , buf_N159_splitterN159ton117n330_1 );
buf_AQFP buf_N165_splitterN165ton129n346_1_( clk_3 , N165 , 0 , buf_N165_splitterN165ton129n346_1 );
buf_AQFP buf_N165_splitterN165ton129n346_2_( clk_5 , buf_N165_splitterN165ton129n346_1 , 0 , buf_N165_splitterN165ton129n346_2 );
buf_AQFP buf_N171_splitterN171ton132n361_1_( clk_3 , N171 , 0 , buf_N171_splitterN171ton132n361_1 );
buf_AQFP buf_N171_splitterN171ton132n361_2_( clk_5 , buf_N171_splitterN171ton132n361_1 , 0 , buf_N171_splitterN171ton132n361_2 );
buf_AQFP buf_N171_splitterN171ton132n361_3_( clk_7 , buf_N171_splitterN171ton132n361_2 , 0 , buf_N171_splitterN171ton132n361_3 );
buf_AQFP buf_N177_splitterN177ton117n315_1_( clk_3 , N177 , 0 , buf_N177_splitterN177ton117n315_1 );
buf_AQFP buf_N177_splitterN177ton117n315_2_( clk_4 , buf_N177_splitterN177ton117n315_1 , 0 , buf_N177_splitterN177ton117n315_2 );
buf_AQFP buf_N183_splitterN183ton132n221_1_( clk_3 , N183 , 0 , buf_N183_splitterN183ton132n221_1 );
buf_AQFP buf_N183_splitterN183ton132n221_2_( clk_4 , buf_N183_splitterN183ton132n221_1 , 0 , buf_N183_splitterN183ton132n221_2 );
buf_AQFP buf_N183_splitterN183ton132n221_3_( clk_6 , buf_N183_splitterN183ton132n221_2 , 0 , buf_N183_splitterN183ton132n221_3 );
buf_AQFP buf_N189_splitterN189ton123n236_1_( clk_3 , N189 , 0 , buf_N189_splitterN189ton123n236_1 );
buf_AQFP buf_N195_splitterN195ton123n253_1_( clk_3 , N195 , 0 , buf_N195_splitterN195ton123n253_1 );
buf_AQFP buf_N195_splitterN195ton123n253_2_( clk_4 , buf_N195_splitterN195ton123n253_1 , 0 , buf_N195_splitterN195ton123n253_2 );
buf_AQFP buf_N195_splitterN195ton123n253_3_( clk_5 , buf_N195_splitterN195ton123n253_2 , 0 , buf_N195_splitterN195ton123n253_3 );
buf_AQFP buf_N195_splitterN195ton123n253_4_( clk_7 , buf_N195_splitterN195ton123n253_3 , 0 , buf_N195_splitterN195ton123n253_4 );
buf_AQFP buf_N201_splitterN201ton129n180_1_( clk_3 , N201 , 0 , buf_N201_splitterN201ton129n180_1 );
buf_AQFP buf_N207_splitterfromN207_1_( clk_3 , N207 , 0 , buf_N207_splitterfromN207_1 );
buf_AQFP buf_N207_splitterfromN207_2_( clk_4 , buf_N207_splitterfromN207_1 , 0 , buf_N207_splitterfromN207_2 );
buf_AQFP buf_N207_splitterfromN207_3_( clk_5 , buf_N207_splitterfromN207_2 , 0 , buf_N207_splitterfromN207_3 );
buf_AQFP buf_N207_splitterfromN207_4_( clk_6 , buf_N207_splitterfromN207_3 , 0 , buf_N207_splitterfromN207_4 );
buf_AQFP buf_N207_splitterfromN207_5_( clk_7 , buf_N207_splitterfromN207_4 , 0 , buf_N207_splitterfromN207_5 );
buf_AQFP buf_N207_splitterfromN207_6_( clk_1 , buf_N207_splitterfromN207_5 , 0 , buf_N207_splitterfromN207_6 );
buf_AQFP buf_N210_splitterN210ton182n360_1_( clk_3 , N210 , 0 , buf_N210_splitterN210ton182n360_1 );
buf_AQFP buf_N219_splitterN219ton171n355_1_( clk_3 , N219 , 0 , buf_N219_splitterN219ton171n355_1 );
buf_AQFP buf_N219_splitterN219ton171n355_2_( clk_5 , buf_N219_splitterN219ton171n355_1 , 0 , buf_N219_splitterN219ton171n355_2 );
buf_AQFP buf_N219_splitterN219ton171n355_3_( clk_7 , buf_N219_splitterN219ton171n355_2 , 0 , buf_N219_splitterN219ton171n355_3 );
buf_AQFP buf_N219_splitterN219ton171n355_4_( clk_1 , buf_N219_splitterN219ton171n355_3 , 0 , buf_N219_splitterN219ton171n355_4 );
buf_AQFP buf_N219_splitterN219ton171n355_5_( clk_3 , buf_N219_splitterN219ton171n355_4 , 0 , buf_N219_splitterN219ton171n355_5 );
buf_AQFP buf_N228_splitterN228ton173n357_1_( clk_3 , N228 , 0 , buf_N228_splitterN228ton173n357_1 );
buf_AQFP buf_N228_splitterN228ton173n357_2_( clk_5 , buf_N228_splitterN228ton173n357_1 , 0 , buf_N228_splitterN228ton173n357_2 );
buf_AQFP buf_N228_splitterN228ton173n357_3_( clk_7 , buf_N228_splitterN228ton173n357_2 , 0 , buf_N228_splitterN228ton173n357_3 );
buf_AQFP buf_N228_splitterN228ton173n357_4_( clk_1 , buf_N228_splitterN228ton173n357_3 , 0 , buf_N228_splitterN228ton173n357_4 );
buf_AQFP buf_N228_splitterN228ton173n357_5_( clk_3 , buf_N228_splitterN228ton173n357_4 , 0 , buf_N228_splitterN228ton173n357_5 );
buf_AQFP buf_N228_splitterN228ton173n357_6_( clk_4 , buf_N228_splitterN228ton173n357_5 , 0 , buf_N228_splitterN228ton173n357_6 );
buf_AQFP buf_N228_splitterN228ton173n357_7_( clk_5 , buf_N228_splitterN228ton173n357_6 , 0 , buf_N228_splitterN228ton173n357_7 );
buf_AQFP buf_N228_splitterN228ton173n357_8_( clk_6 , buf_N228_splitterN228ton173n357_7 , 0 , buf_N228_splitterN228ton173n357_8 );
buf_AQFP buf_N237_splitterN237ton174n358_1_( clk_3 , N237 , 0 , buf_N237_splitterN237ton174n358_1 );
buf_AQFP buf_N246_splitterN246ton175n359_1_( clk_3 , N246 , 0 , buf_N246_splitterN246ton175n359_1 );
buf_AQFP buf_N246_splitterN246ton175n359_2_( clk_4 , buf_N246_splitterN246ton175n359_1 , 0 , buf_N246_splitterN246ton175n359_2 );
buf_AQFP buf_N246_splitterN246ton175n359_3_( clk_6 , buf_N246_splitterN246ton175n359_2 , 0 , buf_N246_splitterN246ton175n359_3 );
buf_AQFP buf_N246_splitterN246ton175n359_4_( clk_8 , buf_N246_splitterN246ton175n359_3 , 0 , buf_N246_splitterN246ton175n359_4 );
buf_AQFP buf_N246_splitterN246ton175n359_5_( clk_2 , buf_N246_splitterN246ton175n359_4 , 0 , buf_N246_splitterN246ton175n359_5 );
buf_AQFP buf_N255_splitterN255ton181n254_1_( clk_3 , N255 , 0 , buf_N255_splitterN255ton181n254_1 );
buf_AQFP buf_N259_n238_1_( clk_3 , N259 , 0 , buf_N259_n238_1 );
buf_AQFP buf_N259_n238_2_( clk_4 , buf_N259_n238_1 , 0 , buf_N259_n238_2 );
buf_AQFP buf_N260_n254_1_( clk_3 , N260 , 0 , buf_N260_n254_1 );
buf_AQFP buf_N260_n254_2_( clk_5 , buf_N260_n254_1 , 0 , buf_N260_n254_2 );
buf_AQFP buf_N261_splitterN261ton169n201_1_( clk_3 , N261 , 0 , buf_N261_splitterN261ton169n201_1 );
buf_AQFP buf_N261_splitterN261ton169n201_2_( clk_5 , buf_N261_splitterN261ton169n201_1 , 0 , buf_N261_splitterN261ton169n201_2 );
buf_AQFP buf_N261_splitterN261ton169n201_3_( clk_7 , buf_N261_splitterN261ton169n201_2 , 0 , buf_N261_splitterN261ton169n201_3 );
buf_AQFP buf_N261_splitterN261ton169n201_4_( clk_1 , buf_N261_splitterN261ton169n201_3 , 0 , buf_N261_splitterN261ton169n201_4 );
buf_AQFP buf_N267_n181_1_( clk_3 , N267 , 0 , buf_N267_n181_1 );
buf_AQFP buf_N267_n181_2_( clk_5 , buf_N267_n181_1 , 0 , buf_N267_n181_2 );
buf_AQFP buf_N268_splitterN268ton152n331_1_( clk_3 , N268 , 0 , buf_N268_splitterN268ton152n331_1 );
buf_AQFP buf_N51_splitterN51ton159n81_1_( clk_2 , N51 , 0 , buf_N51_splitterN51ton159n81_1 );
buf_AQFP buf_N55_splitterN55ton151n82_1_( clk_2 , N55 , 0 , buf_N55_splitterN55ton151n82_1 );
buf_AQFP buf_N55_splitterN55ton151n82_2_( clk_3 , buf_N55_splitterN55ton151n82_1 , 0 , buf_N55_splitterN55ton151n82_2 );
buf_AQFP buf_N72_n176_1_( clk_3 , N72 , 0 , buf_N72_n176_1 );
buf_AQFP buf_N72_n176_2_( clk_5 , buf_N72_n176_1 , 0 , buf_N72_n176_2 );
buf_AQFP buf_N73_n177_1_( clk_3 , N73 , 0 , buf_N73_n177_1 );
buf_AQFP buf_N73_n177_2_( clk_5 , buf_N73_n177_1 , 0 , buf_N73_n177_2 );
buf_AQFP buf_N74_n87_1_( clk_3 , N74 , 0 , buf_N74_n87_1 );
buf_AQFP buf_N74_n87_2_( clk_5 , buf_N74_n87_1 , 0 , buf_N74_n87_2 );
buf_AQFP buf_N74_n87_3_( clk_7 , buf_N74_n87_2 , 0 , buf_N74_n87_3 );
buf_AQFP buf_N80_splitterN80ton149n76_1_( clk_2 , N80 , 0 , buf_N80_splitterN80ton149n76_1 );
buf_AQFP buf_N80_splitterN80ton149n76_2_( clk_3 , buf_N80_splitterN80ton149n76_1 , 0 , buf_N80_splitterN80ton149n76_2 );
buf_AQFP buf_N89_n89_1_( clk_3 , N89 , 0 , buf_N89_n89_1 );
buf_AQFP buf_N89_n89_2_( clk_5 , buf_N89_n89_1 , 0 , buf_N89_n89_2 );
buf_AQFP buf_N90_n79_1_( clk_3 , N90 , 0 , buf_N90_n79_1 );
buf_AQFP buf_N90_n79_2_( clk_5 , buf_N90_n79_1 , 0 , buf_N90_n79_2 );
buf_AQFP buf_N90_n79_3_( clk_7 , buf_N90_n79_2 , 0 , buf_N90_n79_3 );
buf_AQFP buf_N90_n79_4_( clk_1 , buf_N90_n79_3 , 0 , buf_N90_n79_4 );
buf_AQFP buf_N91_splitterN91ton262n94_1_( clk_3 , N91 , 0 , buf_N91_splitterN91ton262n94_1 );
buf_AQFP buf_N91_splitterN91ton262n94_2_( clk_5 , buf_N91_splitterN91ton262n94_1 , 0 , buf_N91_splitterN91ton262n94_2 );
buf_AQFP buf_n62_N388_1_( clk_3 , n62 , 0 , buf_n62_N388_1 );
buf_AQFP buf_n62_N388_2_( clk_5 , buf_n62_N388_1 , 0 , buf_n62_N388_2 );
buf_AQFP buf_n62_N388_3_( clk_7 , buf_n62_N388_2 , 0 , buf_n62_N388_3 );
buf_AQFP buf_n62_N388_4_( clk_1 , buf_n62_N388_3 , 0 , buf_n62_N388_4 );
buf_AQFP buf_n62_N388_5_( clk_3 , buf_n62_N388_4 , 0 , buf_n62_N388_5 );
buf_AQFP buf_n62_N388_6_( clk_5 , buf_n62_N388_5 , 0 , buf_n62_N388_6 );
buf_AQFP buf_n62_N388_7_( clk_7 , buf_n62_N388_6 , 0 , buf_n62_N388_7 );
buf_AQFP buf_n62_N388_8_( clk_1 , buf_n62_N388_7 , 0 , buf_n62_N388_8 );
buf_AQFP buf_n62_N388_9_( clk_3 , buf_n62_N388_8 , 0 , buf_n62_N388_9 );
buf_AQFP buf_n62_N388_10_( clk_5 , buf_n62_N388_9 , 0 , buf_n62_N388_10 );
buf_AQFP buf_n62_N388_11_( clk_7 , buf_n62_N388_10 , 0 , buf_n62_N388_11 );
buf_AQFP buf_n62_N388_12_( clk_1 , buf_n62_N388_11 , 0 , buf_n62_N388_12 );
buf_AQFP buf_n62_N388_13_( clk_3 , buf_n62_N388_12 , 0 , buf_n62_N388_13 );
buf_AQFP buf_n62_N388_14_( clk_5 , buf_n62_N388_13 , 0 , buf_n62_N388_14 );
buf_AQFP buf_n62_N388_15_( clk_7 , buf_n62_N388_14 , 0 , buf_n62_N388_15 );
buf_AQFP buf_n62_N388_16_( clk_1 , buf_n62_N388_15 , 0 , buf_n62_N388_16 );
buf_AQFP buf_n62_N388_17_( clk_3 , buf_n62_N388_16 , 0 , buf_n62_N388_17 );
buf_AQFP buf_n62_N388_18_( clk_4 , buf_n62_N388_17 , 0 , buf_n62_N388_18 );
buf_AQFP buf_n63_splitterfromn63_1_( clk_5 , n63 , 0 , buf_n63_splitterfromn63_1 );
buf_AQFP buf_n63_splitterfromn63_2_( clk_7 , buf_n63_splitterfromn63_1 , 0 , buf_n63_splitterfromn63_2 );
buf_AQFP buf_n64_N389_1_( clk_2 , n64 , 0 , buf_n64_N389_1 );
buf_AQFP buf_n64_N389_2_( clk_4 , buf_n64_N389_1 , 0 , buf_n64_N389_2 );
buf_AQFP buf_n64_N389_3_( clk_6 , buf_n64_N389_2 , 0 , buf_n64_N389_3 );
buf_AQFP buf_n64_N389_4_( clk_8 , buf_n64_N389_3 , 0 , buf_n64_N389_4 );
buf_AQFP buf_n64_N389_5_( clk_2 , buf_n64_N389_4 , 0 , buf_n64_N389_5 );
buf_AQFP buf_n64_N389_6_( clk_4 , buf_n64_N389_5 , 0 , buf_n64_N389_6 );
buf_AQFP buf_n64_N389_7_( clk_6 , buf_n64_N389_6 , 0 , buf_n64_N389_7 );
buf_AQFP buf_n64_N389_8_( clk_8 , buf_n64_N389_7 , 0 , buf_n64_N389_8 );
buf_AQFP buf_n64_N389_9_( clk_2 , buf_n64_N389_8 , 0 , buf_n64_N389_9 );
buf_AQFP buf_n64_N389_10_( clk_4 , buf_n64_N389_9 , 0 , buf_n64_N389_10 );
buf_AQFP buf_n64_N389_11_( clk_6 , buf_n64_N389_10 , 0 , buf_n64_N389_11 );
buf_AQFP buf_n64_N389_12_( clk_8 , buf_n64_N389_11 , 0 , buf_n64_N389_12 );
buf_AQFP buf_n64_N389_13_( clk_2 , buf_n64_N389_12 , 0 , buf_n64_N389_13 );
buf_AQFP buf_n64_N389_14_( clk_4 , buf_n64_N389_13 , 0 , buf_n64_N389_14 );
buf_AQFP buf_n64_N389_15_( clk_6 , buf_n64_N389_14 , 0 , buf_n64_N389_15 );
buf_AQFP buf_n64_N389_16_( clk_8 , buf_n64_N389_15 , 0 , buf_n64_N389_16 );
buf_AQFP buf_n64_N389_17_( clk_2 , buf_n64_N389_16 , 0 , buf_n64_N389_17 );
buf_AQFP buf_n64_N389_18_( clk_4 , buf_n64_N389_17 , 0 , buf_n64_N389_18 );
buf_AQFP buf_n65_splittern65toN390n80_1_( clk_4 , n65 , 0 , buf_n65_splittern65toN390n80_1 );
buf_AQFP buf_n65_splittern65toN390n80_2_( clk_6 , buf_n65_splittern65toN390n80_1 , 0 , buf_n65_splittern65toN390n80_2 );
buf_AQFP buf_n65_splittern65toN390n80_3_( clk_8 , buf_n65_splittern65toN390n80_2 , 0 , buf_n65_splittern65toN390n80_3 );
buf_AQFP buf_n65_splittern65toN390n80_4_( clk_2 , buf_n65_splittern65toN390n80_3 , 0 , buf_n65_splittern65toN390n80_4 );
buf_AQFP buf_n65_splittern65toN390n80_5_( clk_4 , buf_n65_splittern65toN390n80_4 , 0 , buf_n65_splittern65toN390n80_5 );
buf_AQFP buf_n65_splittern65toN390n80_6_( clk_6 , buf_n65_splittern65toN390n80_5 , 0 , buf_n65_splittern65toN390n80_6 );
buf_AQFP buf_n65_splittern65toN390n80_7_( clk_8 , buf_n65_splittern65toN390n80_6 , 0 , buf_n65_splittern65toN390n80_7 );
buf_AQFP buf_n65_splittern65toN390n80_8_( clk_2 , buf_n65_splittern65toN390n80_7 , 0 , buf_n65_splittern65toN390n80_8 );
buf_AQFP buf_n65_splittern65toN390n80_9_( clk_4 , buf_n65_splittern65toN390n80_8 , 0 , buf_n65_splittern65toN390n80_9 );
buf_AQFP buf_n65_splittern65toN390n80_10_( clk_6 , buf_n65_splittern65toN390n80_9 , 0 , buf_n65_splittern65toN390n80_10 );
buf_AQFP buf_n65_splittern65toN390n80_11_( clk_8 , buf_n65_splittern65toN390n80_10 , 0 , buf_n65_splittern65toN390n80_11 );
buf_AQFP buf_n65_splittern65toN390n80_12_( clk_2 , buf_n65_splittern65toN390n80_11 , 0 , buf_n65_splittern65toN390n80_12 );
buf_AQFP buf_n65_splittern65toN390n80_13_( clk_4 , buf_n65_splittern65toN390n80_12 , 0 , buf_n65_splittern65toN390n80_13 );
buf_AQFP buf_n65_splittern65toN390n80_14_( clk_6 , buf_n65_splittern65toN390n80_13 , 0 , buf_n65_splittern65toN390n80_14 );
buf_AQFP buf_n65_splittern65toN390n80_15_( clk_8 , buf_n65_splittern65toN390n80_14 , 0 , buf_n65_splittern65toN390n80_15 );
buf_AQFP buf_n66_N391_1_( clk_5 , n66 , 0 , buf_n66_N391_1 );
buf_AQFP buf_n66_N391_2_( clk_7 , buf_n66_N391_1 , 0 , buf_n66_N391_2 );
buf_AQFP buf_n66_N391_3_( clk_8 , buf_n66_N391_2 , 0 , buf_n66_N391_3 );
buf_AQFP buf_n66_N391_4_( clk_2 , buf_n66_N391_3 , 0 , buf_n66_N391_4 );
buf_AQFP buf_n66_N391_5_( clk_4 , buf_n66_N391_4 , 0 , buf_n66_N391_5 );
buf_AQFP buf_n66_N391_6_( clk_6 , buf_n66_N391_5 , 0 , buf_n66_N391_6 );
buf_AQFP buf_n66_N391_7_( clk_8 , buf_n66_N391_6 , 0 , buf_n66_N391_7 );
buf_AQFP buf_n66_N391_8_( clk_2 , buf_n66_N391_7 , 0 , buf_n66_N391_8 );
buf_AQFP buf_n66_N391_9_( clk_4 , buf_n66_N391_8 , 0 , buf_n66_N391_9 );
buf_AQFP buf_n66_N391_10_( clk_6 , buf_n66_N391_9 , 0 , buf_n66_N391_10 );
buf_AQFP buf_n66_N391_11_( clk_8 , buf_n66_N391_10 , 0 , buf_n66_N391_11 );
buf_AQFP buf_n66_N391_12_( clk_2 , buf_n66_N391_11 , 0 , buf_n66_N391_12 );
buf_AQFP buf_n66_N391_13_( clk_4 , buf_n66_N391_12 , 0 , buf_n66_N391_13 );
buf_AQFP buf_n66_N391_14_( clk_6 , buf_n66_N391_13 , 0 , buf_n66_N391_14 );
buf_AQFP buf_n66_N391_15_( clk_8 , buf_n66_N391_14 , 0 , buf_n66_N391_15 );
buf_AQFP buf_n66_N391_16_( clk_2 , buf_n66_N391_15 , 0 , buf_n66_N391_16 );
buf_AQFP buf_n66_N391_17_( clk_4 , buf_n66_N391_16 , 0 , buf_n66_N391_17 );
buf_AQFP buf_n66_N391_18_( clk_6 , buf_n66_N391_17 , 0 , buf_n66_N391_18 );
buf_AQFP buf_n66_N391_19_( clk_8 , buf_n66_N391_18 , 0 , buf_n66_N391_19 );
buf_AQFP buf_n66_N391_20_( clk_2 , buf_n66_N391_19 , 0 , buf_n66_N391_20 );
buf_AQFP buf_n66_N391_21_( clk_4 , buf_n66_N391_20 , 0 , buf_n66_N391_21 );
buf_AQFP buf_n67_splittern67ton160n83_1_( clk_4 , n67 , 0 , buf_n67_splittern67ton160n83_1 );
buf_AQFP buf_n68_splitterfromn68_1_( clk_1 , n68 , 0 , buf_n68_splitterfromn68_1 );
buf_AQFP buf_n68_splitterfromn68_2_( clk_3 , buf_n68_splitterfromn68_1 , 0 , buf_n68_splitterfromn68_2 );
buf_AQFP buf_n68_splitterfromn68_3_( clk_5 , buf_n68_splitterfromn68_2 , 0 , buf_n68_splitterfromn68_3 );
buf_AQFP buf_n68_splitterfromn68_4_( clk_7 , buf_n68_splitterfromn68_3 , 0 , buf_n68_splitterfromn68_4 );
buf_AQFP buf_n69_N418_1_( clk_7 , n69 , 0 , buf_n69_N418_1 );
buf_AQFP buf_n69_N418_2_( clk_1 , buf_n69_N418_1 , 0 , buf_n69_N418_2 );
buf_AQFP buf_n69_N418_3_( clk_3 , buf_n69_N418_2 , 0 , buf_n69_N418_3 );
buf_AQFP buf_n69_N418_4_( clk_5 , buf_n69_N418_3 , 0 , buf_n69_N418_4 );
buf_AQFP buf_n69_N418_5_( clk_7 , buf_n69_N418_4 , 0 , buf_n69_N418_5 );
buf_AQFP buf_n69_N418_6_( clk_1 , buf_n69_N418_5 , 0 , buf_n69_N418_6 );
buf_AQFP buf_n69_N418_7_( clk_3 , buf_n69_N418_6 , 0 , buf_n69_N418_7 );
buf_AQFP buf_n71_splitterfromn71_1_( clk_5 , n71 , 0 , buf_n71_splitterfromn71_1 );
buf_AQFP buf_n71_splitterfromn71_2_( clk_7 , buf_n71_splitterfromn71_1 , 0 , buf_n71_splitterfromn71_2 );
buf_AQFP buf_n71_splitterfromn71_3_( clk_1 , buf_n71_splitterfromn71_2 , 0 , buf_n71_splitterfromn71_3 );
buf_AQFP buf_n71_splitterfromn71_4_( clk_3 , buf_n71_splitterfromn71_3 , 0 , buf_n71_splitterfromn71_4 );
buf_AQFP buf_n71_splitterfromn71_5_( clk_5 , buf_n71_splitterfromn71_4 , 0 , buf_n71_splitterfromn71_5 );
buf_AQFP buf_n72_N419_1_( clk_4 , n72 , 0 , buf_n72_N419_1 );
buf_AQFP buf_n73_splitterfromn73_1_( clk_4 , n73 , 0 , buf_n73_splitterfromn73_1 );
buf_AQFP buf_n74_N420_1_( clk_1 , n74 , 0 , buf_n74_N420_1 );
buf_AQFP buf_n74_N420_2_( clk_3 , buf_n74_N420_1 , 0 , buf_n74_N420_2 );
buf_AQFP buf_n74_N420_3_( clk_5 , buf_n74_N420_2 , 0 , buf_n74_N420_3 );
buf_AQFP buf_n74_N420_4_( clk_7 , buf_n74_N420_3 , 0 , buf_n74_N420_4 );
buf_AQFP buf_n74_N420_5_( clk_1 , buf_n74_N420_4 , 0 , buf_n74_N420_5 );
buf_AQFP buf_n74_N420_6_( clk_3 , buf_n74_N420_5 , 0 , buf_n74_N420_6 );
buf_AQFP buf_n74_N420_7_( clk_5 , buf_n74_N420_6 , 0 , buf_n74_N420_7 );
buf_AQFP buf_n74_N420_8_( clk_7 , buf_n74_N420_7 , 0 , buf_n74_N420_8 );
buf_AQFP buf_n74_N420_9_( clk_1 , buf_n74_N420_8 , 0 , buf_n74_N420_9 );
buf_AQFP buf_n74_N420_10_( clk_3 , buf_n74_N420_9 , 0 , buf_n74_N420_10 );
buf_AQFP buf_n74_N420_11_( clk_5 , buf_n74_N420_10 , 0 , buf_n74_N420_11 );
buf_AQFP buf_n74_N420_12_( clk_7 , buf_n74_N420_11 , 0 , buf_n74_N420_12 );
buf_AQFP buf_n74_N420_13_( clk_1 , buf_n74_N420_12 , 0 , buf_n74_N420_13 );
buf_AQFP buf_n74_N420_14_( clk_3 , buf_n74_N420_13 , 0 , buf_n74_N420_14 );
buf_AQFP buf_n74_N420_15_( clk_5 , buf_n74_N420_14 , 0 , buf_n74_N420_15 );
buf_AQFP buf_n74_N420_16_( clk_7 , buf_n74_N420_15 , 0 , buf_n74_N420_16 );
buf_AQFP buf_n74_N420_17_( clk_1 , buf_n74_N420_16 , 0 , buf_n74_N420_17 );
buf_AQFP buf_n74_N420_18_( clk_3 , buf_n74_N420_17 , 0 , buf_n74_N420_18 );
buf_AQFP buf_n76_N421_1_( clk_1 , n76 , 0 , buf_n76_N421_1 );
buf_AQFP buf_n76_N421_2_( clk_3 , buf_n76_N421_1 , 0 , buf_n76_N421_2 );
buf_AQFP buf_n76_N421_3_( clk_5 , buf_n76_N421_2 , 0 , buf_n76_N421_3 );
buf_AQFP buf_n76_N421_4_( clk_7 , buf_n76_N421_3 , 0 , buf_n76_N421_4 );
buf_AQFP buf_n76_N421_5_( clk_8 , buf_n76_N421_4 , 0 , buf_n76_N421_5 );
buf_AQFP buf_n76_N421_6_( clk_1 , buf_n76_N421_5 , 0 , buf_n76_N421_6 );
buf_AQFP buf_n76_N421_7_( clk_2 , buf_n76_N421_6 , 0 , buf_n76_N421_7 );
buf_AQFP buf_n76_N421_8_( clk_3 , buf_n76_N421_7 , 0 , buf_n76_N421_8 );
buf_AQFP buf_n76_N421_9_( clk_4 , buf_n76_N421_8 , 0 , buf_n76_N421_9 );
buf_AQFP buf_n77_N422_1_( clk_7 , n77 , 0 , buf_n77_N422_1 );
buf_AQFP buf_n77_N422_2_( clk_8 , buf_n77_N422_1 , 0 , buf_n77_N422_2 );
buf_AQFP buf_n77_N422_3_( clk_1 , buf_n77_N422_2 , 0 , buf_n77_N422_3 );
buf_AQFP buf_n77_N422_4_( clk_2 , buf_n77_N422_3 , 0 , buf_n77_N422_4 );
buf_AQFP buf_n77_N422_5_( clk_3 , buf_n77_N422_4 , 0 , buf_n77_N422_5 );
buf_AQFP buf_n77_N422_6_( clk_4 , buf_n77_N422_5 , 0 , buf_n77_N422_6 );
buf_AQFP buf_n77_N422_7_( clk_5 , buf_n77_N422_6 , 0 , buf_n77_N422_7 );
buf_AQFP buf_n77_N422_8_( clk_6 , buf_n77_N422_7 , 0 , buf_n77_N422_8 );
buf_AQFP buf_n77_N422_9_( clk_7 , buf_n77_N422_8 , 0 , buf_n77_N422_9 );
buf_AQFP buf_n77_N422_10_( clk_1 , buf_n77_N422_9 , 0 , buf_n77_N422_10 );
buf_AQFP buf_n77_N422_11_( clk_3 , buf_n77_N422_10 , 0 , buf_n77_N422_11 );
buf_AQFP buf_n77_N422_12_( clk_5 , buf_n77_N422_11 , 0 , buf_n77_N422_12 );
buf_AQFP buf_n77_N422_13_( clk_7 , buf_n77_N422_12 , 0 , buf_n77_N422_13 );
buf_AQFP buf_n77_N422_14_( clk_1 , buf_n77_N422_13 , 0 , buf_n77_N422_14 );
buf_AQFP buf_n77_N422_15_( clk_3 , buf_n77_N422_14 , 0 , buf_n77_N422_15 );
buf_AQFP buf_n77_N422_16_( clk_5 , buf_n77_N422_15 , 0 , buf_n77_N422_16 );
buf_AQFP buf_n77_N422_17_( clk_6 , buf_n77_N422_16 , 0 , buf_n77_N422_17 );
buf_AQFP buf_n77_N422_18_( clk_8 , buf_n77_N422_17 , 0 , buf_n77_N422_18 );
buf_AQFP buf_n77_N422_19_( clk_2 , buf_n77_N422_18 , 0 , buf_n77_N422_19 );
buf_AQFP buf_n77_N422_20_( clk_4 , buf_n77_N422_19 , 0 , buf_n77_N422_20 );
buf_AQFP buf_n77_N422_21_( clk_6 , buf_n77_N422_20 , 0 , buf_n77_N422_21 );
buf_AQFP buf_n77_N422_22_( clk_8 , buf_n77_N422_21 , 0 , buf_n77_N422_22 );
buf_AQFP buf_n77_N422_23_( clk_2 , buf_n77_N422_22 , 0 , buf_n77_N422_23 );
buf_AQFP buf_n77_N422_24_( clk_4 , buf_n77_N422_23 , 0 , buf_n77_N422_24 );
buf_AQFP buf_n79_N423_1_( clk_4 , n79 , 0 , buf_n79_N423_1 );
buf_AQFP buf_n79_N423_2_( clk_6 , buf_n79_N423_1 , 0 , buf_n79_N423_2 );
buf_AQFP buf_n79_N423_3_( clk_8 , buf_n79_N423_2 , 0 , buf_n79_N423_3 );
buf_AQFP buf_n79_N423_4_( clk_2 , buf_n79_N423_3 , 0 , buf_n79_N423_4 );
buf_AQFP buf_n79_N423_5_( clk_4 , buf_n79_N423_4 , 0 , buf_n79_N423_5 );
buf_AQFP buf_n79_N423_6_( clk_6 , buf_n79_N423_5 , 0 , buf_n79_N423_6 );
buf_AQFP buf_n79_N423_7_( clk_8 , buf_n79_N423_6 , 0 , buf_n79_N423_7 );
buf_AQFP buf_n79_N423_8_( clk_2 , buf_n79_N423_7 , 0 , buf_n79_N423_8 );
buf_AQFP buf_n79_N423_9_( clk_4 , buf_n79_N423_8 , 0 , buf_n79_N423_9 );
buf_AQFP buf_n79_N423_10_( clk_6 , buf_n79_N423_9 , 0 , buf_n79_N423_10 );
buf_AQFP buf_n79_N423_11_( clk_8 , buf_n79_N423_10 , 0 , buf_n79_N423_11 );
buf_AQFP buf_n79_N423_12_( clk_2 , buf_n79_N423_11 , 0 , buf_n79_N423_12 );
buf_AQFP buf_n79_N423_13_( clk_3 , buf_n79_N423_12 , 0 , buf_n79_N423_13 );
buf_AQFP buf_n79_N423_14_( clk_4 , buf_n79_N423_13 , 0 , buf_n79_N423_14 );
buf_AQFP buf_n79_N423_15_( clk_5 , buf_n79_N423_14 , 0 , buf_n79_N423_15 );
buf_AQFP buf_n79_N423_16_( clk_6 , buf_n79_N423_15 , 0 , buf_n79_N423_16 );
buf_AQFP buf_n79_N423_17_( clk_8 , buf_n79_N423_16 , 0 , buf_n79_N423_17 );
buf_AQFP buf_n79_N423_18_( clk_1 , buf_n79_N423_17 , 0 , buf_n79_N423_18 );
buf_AQFP buf_n79_N423_19_( clk_2 , buf_n79_N423_18 , 0 , buf_n79_N423_19 );
buf_AQFP buf_n79_N423_20_( clk_3 , buf_n79_N423_19 , 0 , buf_n79_N423_20 );
buf_AQFP buf_n79_N423_21_( clk_4 , buf_n79_N423_20 , 0 , buf_n79_N423_21 );
buf_AQFP buf_n80_N446_1_( clk_4 , n80 , 0 , buf_n80_N446_1 );
buf_AQFP buf_n84_n85_1_( clk_7 , n84 , 0 , buf_n84_n85_1 );
buf_AQFP buf_n84_n85_2_( clk_1 , buf_n84_n85_1 , 0 , buf_n84_n85_2 );
buf_AQFP buf_n84_n85_3_( clk_3 , buf_n84_n85_2 , 0 , buf_n84_n85_3 );
buf_AQFP buf_n84_n85_4_( clk_5 , buf_n84_n85_3 , 0 , buf_n84_n85_4 );
buf_AQFP buf_n84_n85_5_( clk_7 , buf_n84_n85_4 , 0 , buf_n84_n85_5 );
buf_AQFP buf_n84_n85_6_( clk_1 , buf_n84_n85_5 , 0 , buf_n84_n85_6 );
buf_AQFP buf_n84_n85_7_( clk_3 , buf_n84_n85_6 , 0 , buf_n84_n85_7 );
buf_AQFP buf_n84_n85_8_( clk_5 , buf_n84_n85_7 , 0 , buf_n84_n85_8 );
buf_AQFP buf_n84_n85_9_( clk_7 , buf_n84_n85_8 , 0 , buf_n84_n85_9 );
buf_AQFP buf_n84_n85_10_( clk_1 , buf_n84_n85_9 , 0 , buf_n84_n85_10 );
buf_AQFP buf_n84_n85_11_( clk_3 , buf_n84_n85_10 , 0 , buf_n84_n85_11 );
buf_AQFP buf_n84_n85_12_( clk_5 , buf_n84_n85_11 , 0 , buf_n84_n85_12 );
buf_AQFP buf_n84_n85_13_( clk_7 , buf_n84_n85_12 , 0 , buf_n84_n85_13 );
buf_AQFP buf_n84_n85_14_( clk_1 , buf_n84_n85_13 , 0 , buf_n84_n85_14 );
buf_AQFP buf_n84_n85_15_( clk_3 , buf_n84_n85_14 , 0 , buf_n84_n85_15 );
buf_AQFP buf_n84_n85_16_( clk_5 , buf_n84_n85_15 , 0 , buf_n84_n85_16 );
buf_AQFP buf_n85_N448_1_( clk_8 , n85 , 0 , buf_n85_N448_1 );
buf_AQFP buf_n85_N448_2_( clk_2 , buf_n85_N448_1 , 0 , buf_n85_N448_2 );
buf_AQFP buf_n85_N448_3_( clk_4 , buf_n85_N448_2 , 0 , buf_n85_N448_3 );
buf_AQFP buf_n87_n88_1_( clk_1 , n87 , 0 , buf_n87_n88_1 );
buf_AQFP buf_n88_N449_1_( clk_5 , n88 , 0 , buf_n88_N449_1 );
buf_AQFP buf_n88_N449_2_( clk_7 , buf_n88_N449_1 , 0 , buf_n88_N449_2 );
buf_AQFP buf_n88_N449_3_( clk_1 , buf_n88_N449_2 , 0 , buf_n88_N449_3 );
buf_AQFP buf_n88_N449_4_( clk_3 , buf_n88_N449_3 , 0 , buf_n88_N449_4 );
buf_AQFP buf_n88_N449_5_( clk_5 , buf_n88_N449_4 , 0 , buf_n88_N449_5 );
buf_AQFP buf_n88_N449_6_( clk_7 , buf_n88_N449_5 , 0 , buf_n88_N449_6 );
buf_AQFP buf_n88_N449_7_( clk_1 , buf_n88_N449_6 , 0 , buf_n88_N449_7 );
buf_AQFP buf_n88_N449_8_( clk_3 , buf_n88_N449_7 , 0 , buf_n88_N449_8 );
buf_AQFP buf_n88_N449_9_( clk_5 , buf_n88_N449_8 , 0 , buf_n88_N449_9 );
buf_AQFP buf_n88_N449_10_( clk_7 , buf_n88_N449_9 , 0 , buf_n88_N449_10 );
buf_AQFP buf_n88_N449_11_( clk_1 , buf_n88_N449_10 , 0 , buf_n88_N449_11 );
buf_AQFP buf_n88_N449_12_( clk_3 , buf_n88_N449_11 , 0 , buf_n88_N449_12 );
buf_AQFP buf_n88_N449_13_( clk_5 , buf_n88_N449_12 , 0 , buf_n88_N449_13 );
buf_AQFP buf_n88_N449_14_( clk_7 , buf_n88_N449_13 , 0 , buf_n88_N449_14 );
buf_AQFP buf_n88_N449_15_( clk_1 , buf_n88_N449_14 , 0 , buf_n88_N449_15 );
buf_AQFP buf_n88_N449_16_( clk_3 , buf_n88_N449_15 , 0 , buf_n88_N449_16 );
buf_AQFP buf_n88_N449_17_( clk_4 , buf_n88_N449_16 , 0 , buf_n88_N449_17 );
buf_AQFP buf_n89_N450_1_( clk_8 , n89 , 0 , buf_n89_N450_1 );
buf_AQFP buf_n89_N450_2_( clk_2 , buf_n89_N450_1 , 0 , buf_n89_N450_2 );
buf_AQFP buf_n89_N450_3_( clk_3 , buf_n89_N450_2 , 0 , buf_n89_N450_3 );
buf_AQFP buf_n89_N450_4_( clk_4 , buf_n89_N450_3 , 0 , buf_n89_N450_4 );
buf_AQFP buf_n89_N450_5_( clk_5 , buf_n89_N450_4 , 0 , buf_n89_N450_5 );
buf_AQFP buf_n89_N450_6_( clk_6 , buf_n89_N450_5 , 0 , buf_n89_N450_6 );
buf_AQFP buf_n89_N450_7_( clk_7 , buf_n89_N450_6 , 0 , buf_n89_N450_7 );
buf_AQFP buf_n89_N450_8_( clk_8 , buf_n89_N450_7 , 0 , buf_n89_N450_8 );
buf_AQFP buf_n89_N450_9_( clk_1 , buf_n89_N450_8 , 0 , buf_n89_N450_9 );
buf_AQFP buf_n89_N450_10_( clk_2 , buf_n89_N450_9 , 0 , buf_n89_N450_10 );
buf_AQFP buf_n89_N450_11_( clk_3 , buf_n89_N450_10 , 0 , buf_n89_N450_11 );
buf_AQFP buf_n89_N450_12_( clk_4 , buf_n89_N450_11 , 0 , buf_n89_N450_12 );
buf_AQFP buf_n89_N450_13_( clk_5 , buf_n89_N450_12 , 0 , buf_n89_N450_13 );
buf_AQFP buf_n89_N450_14_( clk_6 , buf_n89_N450_13 , 0 , buf_n89_N450_14 );
buf_AQFP buf_n89_N450_15_( clk_7 , buf_n89_N450_14 , 0 , buf_n89_N450_15 );
buf_AQFP buf_n89_N450_16_( clk_8 , buf_n89_N450_15 , 0 , buf_n89_N450_16 );
buf_AQFP buf_n89_N450_17_( clk_1 , buf_n89_N450_16 , 0 , buf_n89_N450_17 );
buf_AQFP buf_n89_N450_18_( clk_2 , buf_n89_N450_17 , 0 , buf_n89_N450_18 );
buf_AQFP buf_n89_N450_19_( clk_3 , buf_n89_N450_18 , 0 , buf_n89_N450_19 );
buf_AQFP buf_n89_N450_20_( clk_4 , buf_n89_N450_19 , 0 , buf_n89_N450_20 );
buf_AQFP buf_n89_N450_21_( clk_5 , buf_n89_N450_20 , 0 , buf_n89_N450_21 );
buf_AQFP buf_n89_N450_22_( clk_6 , buf_n89_N450_21 , 0 , buf_n89_N450_22 );
buf_AQFP buf_n89_N450_23_( clk_7 , buf_n89_N450_22 , 0 , buf_n89_N450_23 );
buf_AQFP buf_n89_N450_24_( clk_8 , buf_n89_N450_23 , 0 , buf_n89_N450_24 );
buf_AQFP buf_n89_N450_25_( clk_1 , buf_n89_N450_24 , 0 , buf_n89_N450_25 );
buf_AQFP buf_n89_N450_26_( clk_2 , buf_n89_N450_25 , 0 , buf_n89_N450_26 );
buf_AQFP buf_n89_N450_27_( clk_3 , buf_n89_N450_26 , 0 , buf_n89_N450_27 );
buf_AQFP buf_n89_N450_28_( clk_4 , buf_n89_N450_27 , 0 , buf_n89_N450_28 );
buf_AQFP buf_n89_N450_29_( clk_5 , buf_n89_N450_28 , 0 , buf_n89_N450_29 );
buf_AQFP buf_n89_N450_30_( clk_6 , buf_n89_N450_29 , 0 , buf_n89_N450_30 );
buf_AQFP buf_n89_N450_31_( clk_7 , buf_n89_N450_30 , 0 , buf_n89_N450_31 );
buf_AQFP buf_n89_N450_32_( clk_8 , buf_n89_N450_31 , 0 , buf_n89_N450_32 );
buf_AQFP buf_n89_N450_33_( clk_1 , buf_n89_N450_32 , 0 , buf_n89_N450_33 );
buf_AQFP buf_n89_N450_34_( clk_2 , buf_n89_N450_33 , 0 , buf_n89_N450_34 );
buf_AQFP buf_n89_N450_35_( clk_3 , buf_n89_N450_34 , 0 , buf_n89_N450_35 );
buf_AQFP buf_n89_N450_36_( clk_4 , buf_n89_N450_35 , 0 , buf_n89_N450_36 );
buf_AQFP buf_n93_n95_1_( clk_2 , n93 , 0 , buf_n93_n95_1 );
buf_AQFP buf_n94_n95_1_( clk_2 , n94 , 0 , buf_n94_n95_1 );
buf_AQFP buf_n95_splitterfromn95_1_( clk_6 , n95 , 0 , buf_n95_splitterfromn95_1 );
buf_AQFP buf_n95_splitterfromn95_2_( clk_8 , buf_n95_splitterfromn95_1 , 0 , buf_n95_splitterfromn95_2 );
buf_AQFP buf_n95_splitterfromn95_3_( clk_2 , buf_n95_splitterfromn95_2 , 0 , buf_n95_splitterfromn95_3 );
buf_AQFP buf_n113_splitterfromn113_1_( clk_2 , n113 , 0 , buf_n113_splitterfromn113_1 );
buf_AQFP buf_n113_splitterfromn113_2_( clk_4 , buf_n113_splitterfromn113_1 , 0 , buf_n113_splitterfromn113_2 );
buf_AQFP buf_n115_n116_1_( clk_2 , n115 , 0 , buf_n115_n116_1 );
buf_AQFP buf_n115_n116_2_( clk_4 , buf_n115_n116_1 , 0 , buf_n115_n116_2 );
buf_AQFP buf_n115_n116_3_( clk_6 , buf_n115_n116_2 , 0 , buf_n115_n116_3 );
buf_AQFP buf_n115_n116_4_( clk_8 , buf_n115_n116_3 , 0 , buf_n115_n116_4 );
buf_AQFP buf_n116_N767_1_( clk_4 , n116 , 0 , buf_n116_N767_1 );
buf_AQFP buf_n119_splitterfromn119_1_( clk_1 , n119 , 0 , buf_n119_splitterfromn119_1 );
buf_AQFP buf_n122_splitterfromn122_1_( clk_8 , n122 , 0 , buf_n122_splitterfromn122_1 );
buf_AQFP buf_n122_splitterfromn122_2_( clk_2 , buf_n122_splitterfromn122_1 , 0 , buf_n122_splitterfromn122_2 );
buf_AQFP buf_n122_splitterfromn122_3_( clk_4 , buf_n122_splitterfromn122_2 , 0 , buf_n122_splitterfromn122_3 );
buf_AQFP buf_n140_splitterfromn140_1_( clk_6 , n140 , 0 , buf_n140_splitterfromn140_1 );
buf_AQFP buf_n140_splitterfromn140_2_( clk_7 , buf_n140_splitterfromn140_1 , 0 , buf_n140_splitterfromn140_2 );
buf_AQFP buf_n143_N768_1_( clk_5 , n143 , 0 , buf_n143_N768_1 );
buf_AQFP buf_n143_N768_2_( clk_7 , buf_n143_N768_1 , 0 , buf_n143_N768_2 );
buf_AQFP buf_n143_N768_3_( clk_1 , buf_n143_N768_2 , 0 , buf_n143_N768_3 );
buf_AQFP buf_n143_N768_4_( clk_2 , buf_n143_N768_3 , 0 , buf_n143_N768_4 );
buf_AQFP buf_n143_N768_5_( clk_4 , buf_n143_N768_4 , 0 , buf_n143_N768_5 );
buf_AQFP buf_n143_N768_6_( clk_5 , buf_n143_N768_5 , 0 , buf_n143_N768_6 );
buf_AQFP buf_n143_N768_7_( clk_7 , buf_n143_N768_6 , 0 , buf_n143_N768_7 );
buf_AQFP buf_n143_N768_8_( clk_8 , buf_n143_N768_7 , 0 , buf_n143_N768_8 );
buf_AQFP buf_n143_N768_9_( clk_2 , buf_n143_N768_8 , 0 , buf_n143_N768_9 );
buf_AQFP buf_n143_N768_10_( clk_4 , buf_n143_N768_9 , 0 , buf_n143_N768_10 );
buf_AQFP buf_n153_n155_1_( clk_6 , n153 , 0 , buf_n153_n155_1 );
buf_AQFP buf_n154_n155_1_( clk_6 , n154 , 0 , buf_n154_n155_1 );
buf_AQFP buf_n181_n183_1_( clk_1 , n181 , 0 , buf_n181_n183_1 );
buf_AQFP buf_n181_n183_2_( clk_2 , buf_n181_n183_1 , 0 , buf_n181_n183_2 );
buf_AQFP buf_n182_n183_1_( clk_1 , n182 , 0 , buf_n182_n183_1 );
buf_AQFP buf_n183_n184_1_( clk_4 , n183 , 0 , buf_n183_n184_1 );
buf_AQFP buf_n184_n185_1_( clk_8 , n184 , 0 , buf_n184_n185_1 );
buf_AQFP buf_n187_n188_1_( clk_5 , n187 , 0 , buf_n187_n188_1 );
buf_AQFP buf_n188_N850_1_( clk_1 , n188 , 0 , buf_n188_N850_1 );
buf_AQFP buf_n188_N850_2_( clk_3 , buf_n188_N850_1 , 0 , buf_n188_N850_2 );
buf_AQFP buf_n188_N850_3_( clk_5 , buf_n188_N850_2 , 0 , buf_n188_N850_3 );
buf_AQFP buf_n188_N850_4_( clk_7 , buf_n188_N850_3 , 0 , buf_n188_N850_4 );
buf_AQFP buf_n188_N850_5_( clk_1 , buf_n188_N850_4 , 0 , buf_n188_N850_5 );
buf_AQFP buf_n188_N850_6_( clk_3 , buf_n188_N850_5 , 0 , buf_n188_N850_6 );
buf_AQFP buf_n188_N850_7_( clk_5 , buf_n188_N850_6 , 0 , buf_n188_N850_7 );
buf_AQFP buf_n188_N850_8_( clk_7 , buf_n188_N850_7 , 0 , buf_n188_N850_8 );
buf_AQFP buf_n188_N850_9_( clk_8 , buf_n188_N850_8 , 0 , buf_n188_N850_9 );
buf_AQFP buf_n188_N850_10_( clk_1 , buf_n188_N850_9 , 0 , buf_n188_N850_10 );
buf_AQFP buf_n188_N850_11_( clk_2 , buf_n188_N850_10 , 0 , buf_n188_N850_11 );
buf_AQFP buf_n188_N850_12_( clk_4 , buf_n188_N850_11 , 0 , buf_n188_N850_12 );
buf_AQFP buf_n217_n227_1_( clk_7 , n217 , 0 , buf_n217_n227_1 );
buf_AQFP buf_n217_n227_2_( clk_1 , buf_n217_n227_1 , 0 , buf_n217_n227_2 );
buf_AQFP buf_n217_n227_3_( clk_2 , buf_n217_n227_2 , 0 , buf_n217_n227_3 );
buf_AQFP buf_n217_n227_4_( clk_4 , buf_n217_n227_3 , 0 , buf_n217_n227_4 );
buf_AQFP buf_n217_n227_5_( clk_5 , buf_n217_n227_4 , 0 , buf_n217_n227_5 );
buf_AQFP buf_n218_n226_1_( clk_6 , n218 , 0 , buf_n218_n226_1 );
buf_AQFP buf_n218_n226_2_( clk_8 , buf_n218_n226_1 , 0 , buf_n218_n226_2 );
buf_AQFP buf_n218_n226_3_( clk_2 , buf_n218_n226_2 , 0 , buf_n218_n226_3 );
buf_AQFP buf_n222_n223_1_( clk_1 , n222 , 0 , buf_n222_n223_1 );
buf_AQFP buf_n222_n223_2_( clk_3 , buf_n222_n223_1 , 0 , buf_n222_n223_2 );
buf_AQFP buf_n222_n223_3_( clk_5 , buf_n222_n223_2 , 0 , buf_n222_n223_3 );
buf_AQFP buf_n223_n224_1_( clk_7 , n223 , 0 , buf_n223_n224_1 );
buf_AQFP buf_n223_n224_2_( clk_8 , buf_n223_n224_1 , 0 , buf_n223_n224_2 );
buf_AQFP buf_n223_n224_3_( clk_1 , buf_n223_n224_2 , 0 , buf_n223_n224_3 );
buf_AQFP buf_n224_n225_1_( clk_3 , n224 , 0 , buf_n224_n225_1 );
buf_AQFP buf_n225_n226_1_( clk_7 , n225 , 0 , buf_n225_n226_1 );
buf_AQFP buf_n225_n226_2_( clk_1 , buf_n225_n226_1 , 0 , buf_n225_n226_2 );
buf_AQFP buf_n226_n227_1_( clk_4 , n226 , 0 , buf_n226_n227_1 );
buf_AQFP buf_n226_n227_2_( clk_6 , buf_n226_n227_1 , 0 , buf_n226_n227_2 );
buf_AQFP buf_n226_n227_3_( clk_8 , buf_n226_n227_2 , 0 , buf_n226_n227_3 );
buf_AQFP buf_n226_n227_4_( clk_2 , buf_n226_n227_3 , 0 , buf_n226_n227_4 );
buf_AQFP buf_n226_n227_5_( clk_4 , buf_n226_n227_4 , 0 , buf_n226_n227_5 );
buf_AQFP buf_n226_n227_6_( clk_5 , buf_n226_n227_5 , 0 , buf_n226_n227_6 );
buf_AQFP buf_n227_N863_1_( clk_7 , n227 , 0 , buf_n227_N863_1 );
buf_AQFP buf_n227_N863_2_( clk_8 , buf_n227_N863_1 , 0 , buf_n227_N863_2 );
buf_AQFP buf_n227_N863_3_( clk_1 , buf_n227_N863_2 , 0 , buf_n227_N863_3 );
buf_AQFP buf_n227_N863_4_( clk_2 , buf_n227_N863_3 , 0 , buf_n227_N863_4 );
buf_AQFP buf_n227_N863_5_( clk_3 , buf_n227_N863_4 , 0 , buf_n227_N863_5 );
buf_AQFP buf_n227_N863_6_( clk_4 , buf_n227_N863_5 , 0 , buf_n227_N863_6 );
buf_AQFP buf_n237_n239_1_( clk_1 , n237 , 0 , buf_n237_n239_1 );
buf_AQFP buf_n238_n239_1_( clk_7 , n238 , 0 , buf_n238_n239_1 );
buf_AQFP buf_n238_n239_2_( clk_8 , buf_n238_n239_1 , 0 , buf_n238_n239_2 );
buf_AQFP buf_n238_n239_3_( clk_1 , buf_n238_n239_2 , 0 , buf_n238_n239_3 );
buf_AQFP buf_n239_n240_1_( clk_3 , n239 , 0 , buf_n239_n240_1 );
buf_AQFP buf_n239_n240_2_( clk_4 , buf_n239_n240_1 , 0 , buf_n239_n240_2 );
buf_AQFP buf_n239_n240_3_( clk_5 , buf_n239_n240_2 , 0 , buf_n239_n240_3 );
buf_AQFP buf_n239_n240_4_( clk_6 , buf_n239_n240_3 , 0 , buf_n239_n240_4 );
buf_AQFP buf_n243_n244_1_( clk_6 , n243 , 0 , buf_n243_n244_1 );
buf_AQFP buf_n243_n244_2_( clk_7 , buf_n243_n244_1 , 0 , buf_n243_n244_2 );
buf_AQFP buf_n243_n244_3_( clk_1 , buf_n243_n244_2 , 0 , buf_n243_n244_3 );
buf_AQFP buf_n244_N864_1_( clk_3 , n244 , 0 , buf_n244_N864_1 );
buf_AQFP buf_n244_N864_2_( clk_4 , buf_n244_N864_1 , 0 , buf_n244_N864_2 );
buf_AQFP buf_n244_N864_3_( clk_5 , buf_n244_N864_2 , 0 , buf_n244_N864_3 );
buf_AQFP buf_n244_N864_4_( clk_6 , buf_n244_N864_3 , 0 , buf_n244_N864_4 );
buf_AQFP buf_n244_N864_5_( clk_7 , buf_n244_N864_4 , 0 , buf_n244_N864_5 );
buf_AQFP buf_n244_N864_6_( clk_8 , buf_n244_N864_5 , 0 , buf_n244_N864_6 );
buf_AQFP buf_n244_N864_7_( clk_1 , buf_n244_N864_6 , 0 , buf_n244_N864_7 );
buf_AQFP buf_n244_N864_8_( clk_2 , buf_n244_N864_7 , 0 , buf_n244_N864_8 );
buf_AQFP buf_n244_N864_9_( clk_3 , buf_n244_N864_8 , 0 , buf_n244_N864_9 );
buf_AQFP buf_n244_N864_10_( clk_4 , buf_n244_N864_9 , 0 , buf_n244_N864_10 );
buf_AQFP buf_n244_N864_11_( clk_5 , buf_n244_N864_10 , 0 , buf_n244_N864_11 );
buf_AQFP buf_n244_N864_12_( clk_6 , buf_n244_N864_11 , 0 , buf_n244_N864_12 );
buf_AQFP buf_n244_N864_13_( clk_8 , buf_n244_N864_12 , 0 , buf_n244_N864_13 );
buf_AQFP buf_n244_N864_14_( clk_2 , buf_n244_N864_13 , 0 , buf_n244_N864_14 );
buf_AQFP buf_n244_N864_15_( clk_4 , buf_n244_N864_14 , 0 , buf_n244_N864_15 );
buf_AQFP buf_n256_n257_1_( clk_2 , n256 , 0 , buf_n256_n257_1 );
buf_AQFP buf_n256_n257_2_( clk_4 , buf_n256_n257_1 , 0 , buf_n256_n257_2 );
buf_AQFP buf_n256_n257_3_( clk_6 , buf_n256_n257_2 , 0 , buf_n256_n257_3 );
buf_AQFP buf_n256_n257_4_( clk_7 , buf_n256_n257_3 , 0 , buf_n256_n257_4 );
buf_AQFP buf_n256_n257_5_( clk_8 , buf_n256_n257_4 , 0 , buf_n256_n257_5 );
buf_AQFP buf_n259_n260_1_( clk_4 , n259 , 0 , buf_n259_n260_1 );
buf_AQFP buf_n261_N865_1_( clk_1 , n261 , 0 , buf_n261_N865_1 );
buf_AQFP buf_n261_N865_2_( clk_3 , buf_n261_N865_1 , 0 , buf_n261_N865_2 );
buf_AQFP buf_n261_N865_3_( clk_5 , buf_n261_N865_2 , 0 , buf_n261_N865_3 );
buf_AQFP buf_n261_N865_4_( clk_7 , buf_n261_N865_3 , 0 , buf_n261_N865_4 );
buf_AQFP buf_n261_N865_5_( clk_1 , buf_n261_N865_4 , 0 , buf_n261_N865_5 );
buf_AQFP buf_n261_N865_6_( clk_3 , buf_n261_N865_5 , 0 , buf_n261_N865_6 );
buf_AQFP buf_n261_N865_7_( clk_5 , buf_n261_N865_6 , 0 , buf_n261_N865_7 );
buf_AQFP buf_n261_N865_8_( clk_7 , buf_n261_N865_7 , 0 , buf_n261_N865_8 );
buf_AQFP buf_n261_N865_9_( clk_1 , buf_n261_N865_8 , 0 , buf_n261_N865_9 );
buf_AQFP buf_n261_N865_10_( clk_3 , buf_n261_N865_9 , 0 , buf_n261_N865_10 );
buf_AQFP buf_n261_N865_11_( clk_4 , buf_n261_N865_10 , 0 , buf_n261_N865_11 );
buf_AQFP buf_n265_n266_1_( clk_7 , n265 , 0 , buf_n265_n266_1 );
buf_AQFP buf_n280_splitterfromn280_1_( clk_2 , n280 , 0 , buf_n280_splitterfromn280_1 );
buf_AQFP buf_n280_splitterfromn280_2_( clk_4 , buf_n280_splitterfromn280_1 , 0 , buf_n280_splitterfromn280_2 );
buf_AQFP buf_n280_splitterfromn280_3_( clk_5 , buf_n280_splitterfromn280_2 , 0 , buf_n280_splitterfromn280_3 );
buf_AQFP buf_n280_splitterfromn280_4_( clk_6 , buf_n280_splitterfromn280_3 , 0 , buf_n280_splitterfromn280_4 );
buf_AQFP buf_n306_N866_1_( clk_2 , n306 , 0 , buf_n306_N866_1 );
buf_AQFP buf_n306_N866_2_( clk_4 , buf_n306_N866_1 , 0 , buf_n306_N866_2 );
buf_AQFP buf_n307_splitterfromn307_1_( clk_6 , n307 , 0 , buf_n307_splitterfromn307_1 );
buf_AQFP buf_n316_n317_1_( clk_2 , n316 , 0 , buf_n316_n317_1 );
buf_AQFP buf_n316_n317_2_( clk_4 , buf_n316_n317_1 , 0 , buf_n316_n317_2 );
buf_AQFP buf_n316_n317_3_( clk_5 , buf_n316_n317_2 , 0 , buf_n316_n317_3 );
buf_AQFP buf_n318_n319_1_( clk_1 , n318 , 0 , buf_n318_n319_1 );
buf_AQFP buf_n319_n320_1_( clk_4 , n319 , 0 , buf_n319_n320_1 );
buf_AQFP buf_n319_n320_2_( clk_5 , buf_n319_n320_1 , 0 , buf_n319_n320_2 );
buf_AQFP buf_n319_n320_3_( clk_6 , buf_n319_n320_2 , 0 , buf_n319_n320_3 );
buf_AQFP buf_n319_n320_4_( clk_7 , buf_n319_n320_3 , 0 , buf_n319_n320_4 );
buf_AQFP buf_n319_n320_5_( clk_8 , buf_n319_n320_4 , 0 , buf_n319_n320_5 );
buf_AQFP buf_n319_n320_6_( clk_2 , buf_n319_n320_5 , 0 , buf_n319_n320_6 );
buf_AQFP buf_n319_n320_7_( clk_4 , buf_n319_n320_6 , 0 , buf_n319_n320_7 );
buf_AQFP buf_n319_n320_8_( clk_6 , buf_n319_n320_7 , 0 , buf_n319_n320_8 );
buf_AQFP buf_n321_N874_1_( clk_4 , n321 , 0 , buf_n321_N874_1 );
buf_AQFP buf_n321_N874_2_( clk_5 , buf_n321_N874_1 , 0 , buf_n321_N874_2 );
buf_AQFP buf_n321_N874_3_( clk_6 , buf_n321_N874_2 , 0 , buf_n321_N874_3 );
buf_AQFP buf_n321_N874_4_( clk_7 , buf_n321_N874_3 , 0 , buf_n321_N874_4 );
buf_AQFP buf_n321_N874_5_( clk_8 , buf_n321_N874_4 , 0 , buf_n321_N874_5 );
buf_AQFP buf_n321_N874_6_( clk_2 , buf_n321_N874_5 , 0 , buf_n321_N874_6 );
buf_AQFP buf_n321_N874_7_( clk_4 , buf_n321_N874_6 , 0 , buf_n321_N874_7 );
buf_AQFP buf_n323_n326_1_( clk_7 , n323 , 0 , buf_n323_n326_1 );
buf_AQFP buf_n327_n335_1_( clk_7 , n327 , 0 , buf_n327_n335_1 );
buf_AQFP buf_n331_n332_1_( clk_2 , n331 , 0 , buf_n331_n332_1 );
buf_AQFP buf_n331_n332_2_( clk_4 , buf_n331_n332_1 , 0 , buf_n331_n332_2 );
buf_AQFP buf_n331_n332_3_( clk_6 , buf_n331_n332_2 , 0 , buf_n331_n332_3 );
buf_AQFP buf_n334_n335_1_( clk_3 , n334 , 0 , buf_n334_n335_1 );
buf_AQFP buf_n334_n335_2_( clk_4 , buf_n334_n335_1 , 0 , buf_n334_n335_2 );
buf_AQFP buf_n334_n335_3_( clk_6 , buf_n334_n335_2 , 0 , buf_n334_n335_3 );
buf_AQFP buf_n334_n335_4_( clk_8 , buf_n334_n335_3 , 0 , buf_n334_n335_4 );
buf_AQFP buf_n335_n336_1_( clk_3 , n335 , 0 , buf_n335_n336_1 );
buf_AQFP buf_n335_n336_2_( clk_4 , buf_n335_n336_1 , 0 , buf_n335_n336_2 );
buf_AQFP buf_n335_n336_3_( clk_6 , buf_n335_n336_2 , 0 , buf_n335_n336_3 );
buf_AQFP buf_n335_n336_4_( clk_7 , buf_n335_n336_3 , 0 , buf_n335_n336_4 );
buf_AQFP buf_n335_n336_5_( clk_8 , buf_n335_n336_4 , 0 , buf_n335_n336_5 );
buf_AQFP buf_n335_n336_6_( clk_1 , buf_n335_n336_5 , 0 , buf_n335_n336_6 );
buf_AQFP buf_n335_n336_7_( clk_2 , buf_n335_n336_6 , 0 , buf_n335_n336_7 );
buf_AQFP buf_n335_n336_8_( clk_3 , buf_n335_n336_7 , 0 , buf_n335_n336_8 );
buf_AQFP buf_n335_n336_9_( clk_5 , buf_n335_n336_8 , 0 , buf_n335_n336_9 );
buf_AQFP buf_n335_n336_10_( clk_6 , buf_n335_n336_9 , 0 , buf_n335_n336_10 );
buf_AQFP buf_n335_n336_11_( clk_7 , buf_n335_n336_10 , 0 , buf_n335_n336_11 );
buf_AQFP buf_n335_n336_12_( clk_1 , buf_n335_n336_11 , 0 , buf_n335_n336_12 );
buf_AQFP buf_n337_splittern337ton338n342_1_( clk_1 , n337 , 0 , buf_n337_splittern337ton338n342_1 );
buf_AQFP buf_n337_splittern337ton338n342_2_( clk_3 , buf_n337_splittern337ton338n342_1 , 0 , buf_n337_splittern337ton338n342_2 );
buf_AQFP buf_n337_splittern337ton338n342_3_( clk_4 , buf_n337_splittern337ton338n342_2 , 0 , buf_n337_splittern337ton338n342_3 );
buf_AQFP buf_n345_n347_1_( clk_3 , n345 , 0 , buf_n345_n347_1 );
buf_AQFP buf_n345_n347_2_( clk_5 , buf_n345_n347_1 , 0 , buf_n345_n347_2 );
buf_AQFP buf_n345_n347_3_( clk_6 , buf_n345_n347_2 , 0 , buf_n345_n347_3 );
buf_AQFP buf_n349_n350_1_( clk_3 , n349 , 0 , buf_n349_n350_1 );
buf_AQFP buf_n349_n350_2_( clk_4 , buf_n349_n350_1 , 0 , buf_n349_n350_2 );
buf_AQFP buf_n349_n350_3_( clk_5 , buf_n349_n350_2 , 0 , buf_n349_n350_3 );
buf_AQFP buf_n349_n350_4_( clk_6 , buf_n349_n350_3 , 0 , buf_n349_n350_4 );
buf_AQFP buf_n349_n350_5_( clk_7 , buf_n349_n350_4 , 0 , buf_n349_n350_5 );
buf_AQFP buf_n349_n350_6_( clk_1 , buf_n349_n350_5 , 0 , buf_n349_n350_6 );
buf_AQFP buf_n349_n350_7_( clk_3 , buf_n349_n350_6 , 0 , buf_n349_n350_7 );
buf_AQFP buf_n349_n350_8_( clk_4 , buf_n349_n350_7 , 0 , buf_n349_n350_8 );
buf_AQFP buf_n349_n350_9_( clk_5 , buf_n349_n350_8 , 0 , buf_n349_n350_9 );
buf_AQFP buf_n349_n350_10_( clk_6 , buf_n349_n350_9 , 0 , buf_n349_n350_10 );
buf_AQFP buf_n349_n350_11_( clk_7 , buf_n349_n350_10 , 0 , buf_n349_n350_11 );
buf_AQFP buf_n349_n350_12_( clk_8 , buf_n349_n350_11 , 0 , buf_n349_n350_12 );
buf_AQFP buf_n350_n351_1_( clk_2 , n350 , 0 , buf_n350_n351_1 );
buf_AQFP buf_n350_n351_2_( clk_3 , buf_n350_n351_1 , 0 , buf_n350_n351_2 );
buf_AQFP buf_n350_n351_3_( clk_4 , buf_n350_n351_2 , 0 , buf_n350_n351_3 );
buf_AQFP buf_n350_n351_4_( clk_5 , buf_n350_n351_3 , 0 , buf_n350_n351_4 );
buf_AQFP buf_n350_n351_5_( clk_6 , buf_n350_n351_4 , 0 , buf_n350_n351_5 );
buf_AQFP buf_n350_n351_6_( clk_7 , buf_n350_n351_5 , 0 , buf_n350_n351_6 );
buf_AQFP buf_n351_N879_1_( clk_2 , n351 , 0 , buf_n351_N879_1 );
buf_AQFP buf_n351_N879_2_( clk_4 , buf_n351_N879_1 , 0 , buf_n351_N879_2 );
buf_AQFP buf_n356_n366_1_( clk_4 , n356 , 0 , buf_n356_n366_1 );
buf_AQFP buf_n356_n366_2_( clk_5 , buf_n356_n366_1 , 0 , buf_n356_n366_2 );
buf_AQFP buf_n356_n366_3_( clk_7 , buf_n356_n366_2 , 0 , buf_n356_n366_3 );
buf_AQFP buf_n360_n362_1_( clk_2 , n360 , 0 , buf_n360_n362_1 );
buf_AQFP buf_n360_n362_2_( clk_3 , buf_n360_n362_1 , 0 , buf_n360_n362_2 );
buf_AQFP buf_n360_n362_3_( clk_4 , buf_n360_n362_2 , 0 , buf_n360_n362_3 );
buf_AQFP buf_n360_n362_4_( clk_5 , buf_n360_n362_3 , 0 , buf_n360_n362_4 );
buf_AQFP buf_n362_n363_1_( clk_7 , n362 , 0 , buf_n362_n363_1 );
buf_AQFP buf_n364_n365_1_( clk_3 , n364 , 0 , buf_n364_n365_1 );
buf_AQFP buf_n364_n365_2_( clk_4 , buf_n364_n365_1 , 0 , buf_n364_n365_2 );
buf_AQFP buf_n364_n365_3_( clk_5 , buf_n364_n365_2 , 0 , buf_n364_n365_3 );
buf_AQFP buf_n364_n365_4_( clk_6 , buf_n364_n365_3 , 0 , buf_n364_n365_4 );
buf_AQFP buf_n364_n365_5_( clk_7 , buf_n364_n365_4 , 0 , buf_n364_n365_5 );
buf_AQFP buf_n365_n366_1_( clk_2 , n365 , 0 , buf_n365_n366_1 );
buf_AQFP buf_n365_n366_2_( clk_4 , buf_n365_n366_1 , 0 , buf_n365_n366_2 );
buf_AQFP buf_n365_n366_3_( clk_6 , buf_n365_n366_2 , 0 , buf_n365_n366_3 );
buf_AQFP buf_n365_n366_4_( clk_7 , buf_n365_n366_3 , 0 , buf_n365_n366_4 );
buf_AQFP buf_n365_n366_5_( clk_8 , buf_n365_n366_4 , 0 , buf_n365_n366_5 );
buf_AQFP buf_n365_n366_6_( clk_1 , buf_n365_n366_5 , 0 , buf_n365_n366_6 );
buf_AQFP buf_n365_n366_7_( clk_2 , buf_n365_n366_6 , 0 , buf_n365_n366_7 );
buf_AQFP buf_n365_n366_8_( clk_3 , buf_n365_n366_7 , 0 , buf_n365_n366_8 );
buf_AQFP buf_n365_n366_9_( clk_4 , buf_n365_n366_8 , 0 , buf_n365_n366_9 );
buf_AQFP buf_n365_n366_10_( clk_5 , buf_n365_n366_9 , 0 , buf_n365_n366_10 );
buf_AQFP buf_n365_n366_11_( clk_7 , buf_n365_n366_10 , 0 , buf_n365_n366_11 );
buf_AQFP buf_n366_N880_1_( clk_3 , n366 , 0 , buf_n366_N880_1 );
buf_AQFP buf_splitterN1ton147n70_n147_1_( clk_4 , splitterN1ton147n70 , 0 , buf_splitterN1ton147n70_n147_1 );
buf_AQFP buf_splitterN1ton147n70_n147_2_( clk_6 , buf_splitterN1ton147n70_n147_1 , 0 , buf_splitterN1ton147n70_n147_2 );
buf_AQFP buf_splitterN1ton147n70_n147_3_( clk_7 , buf_splitterN1ton147n70_n147_2 , 0 , buf_splitterN1ton147n70_n147_3 );
buf_AQFP buf_splitterN1ton147n70_n147_4_( clk_8 , buf_splitterN1ton147n70_n147_3 , 0 , buf_splitterN1ton147n70_n147_4 );
buf_AQFP buf_splitterN101ton102n316_n281_1_( clk_6 , splitterN101ton102n316 , 0 , buf_splitterN101ton102n316_n281_1 );
buf_AQFP buf_splitterN101ton102n316_n281_2_( clk_8 , buf_splitterN101ton102n316_n281_1 , 0 , buf_splitterN101ton102n316_n281_2 );
buf_AQFP buf_splitterN101ton102n316_n281_3_( clk_2 , buf_splitterN101ton102n316_n281_2 , 0 , buf_splitterN101ton102n316_n281_3 );
buf_AQFP buf_splitterN101ton102n316_n316_1_( clk_6 , splitterN101ton102n316 , 0 , buf_splitterN101ton102n316_n316_1 );
buf_AQFP buf_splitterN106ton102n289_n289_1_( clk_7 , splitterN106ton102n289 , 0 , buf_splitterN106ton102n289_n289_1 );
buf_AQFP buf_splitterN106ton102n289_n289_2_( clk_1 , buf_splitterN106ton102n289_n289_1 , 0 , buf_splitterN106ton102n289_n289_2 );
buf_AQFP buf_splitterN106ton102n289_n289_3_( clk_2 , buf_splitterN106ton102n289_n289_2 , 0 , buf_splitterN106ton102n289_n289_3 );
buf_AQFP buf_splitterN111ton105n237_n207_1_( clk_7 , splitterN111ton105n237 , 0 , buf_splitterN111ton105n237_n207_1 );
buf_AQFP buf_splitterN111ton105n237_n207_2_( clk_1 , buf_splitterN111ton105n237_n207_1 , 0 , buf_splitterN111ton105n237_n207_2 );
buf_AQFP buf_splitterN111ton105n237_n207_3_( clk_3 , buf_splitterN111ton105n237_n207_2 , 0 , buf_splitterN111ton105n237_n207_3 );
buf_AQFP buf_splitterN116ton105n255_n190_1_( clk_7 , splitterN116ton105n255 , 0 , buf_splitterN116ton105n255_n190_1 );
buf_AQFP buf_splitterN116ton105n255_n190_2_( clk_1 , buf_splitterN116ton105n255_n190_1 , 0 , buf_splitterN116ton105n255_n190_2 );
buf_AQFP buf_splitterN116ton105n255_n255_1_( clk_6 , splitterN116ton105n255 , 0 , buf_splitterN116ton105n255_n255_1 );
buf_AQFP buf_splitterN121ton182n97_n196_1_( clk_7 , splitterN121ton182n97 , 0 , buf_splitterN121ton182n97_n196_1 );
buf_AQFP buf_splitterN121ton182n97_n196_2_( clk_1 , buf_splitterN121ton182n97_n196_1 , 0 , buf_splitterN121ton182n97_n196_2 );
buf_AQFP buf_splitterN121ton182n97_n196_3_( clk_2 , buf_splitterN121ton182n97_n196_2 , 0 , buf_splitterN121ton182n97_n196_3 );
buf_AQFP buf_splitterN126ton100n99_n163_1_( clk_1 , splitterN126ton100n99 , 0 , buf_splitterN126ton100n99_n163_1 );
buf_AQFP buf_splitterfromN13_n68_1_( clk_6 , splitterfromN13 , 0 , buf_splitterfromN13_n68_1 );
buf_AQFP buf_splitterN130ton120n91_n120_1_( clk_4 , splitterN130ton120n91 , 0 , buf_splitterN130ton120n91_n120_1 );
buf_AQFP buf_splitterN130ton120n91_n120_2_( clk_6 , buf_splitterN130ton120n91_n120_1 , 0 , buf_splitterN130ton120n91_n120_2 );
buf_AQFP buf_splitterN130ton120n91_n120_3_( clk_8 , buf_splitterN130ton120n91_n120_2 , 0 , buf_splitterN130ton120n91_n120_3 );
buf_AQFP buf_splitterN130ton120n91_n120_4_( clk_2 , buf_splitterN130ton120n91_n120_3 , 0 , buf_splitterN130ton120n91_n120_4 );
buf_AQFP buf_splitterN130ton120n91_n121_1_( clk_4 , splitterN130ton120n91 , 0 , buf_splitterN130ton120n91_n121_1 );
buf_AQFP buf_splitterN130ton120n91_n121_2_( clk_6 , buf_splitterN130ton120n91_n121_1 , 0 , buf_splitterN130ton120n91_n121_2 );
buf_AQFP buf_splitterN130ton120n91_n121_3_( clk_8 , buf_splitterN130ton120n91_n121_2 , 0 , buf_splitterN130ton120n91_n121_3 );
buf_AQFP buf_splitterN130ton120n91_n121_4_( clk_2 , buf_splitterN130ton120n91_n121_3 , 0 , buf_splitterN130ton120n91_n121_4 );
buf_AQFP buf_splitterN138ton267n291_n267_1_( clk_8 , splitterN138ton267n291 , 0 , buf_splitterN138ton267n291_n267_1 );
buf_AQFP buf_splitterN138ton267n291_n283_1_( clk_8 , splitterN138ton267n291 , 0 , buf_splitterN138ton267n291_n283_1 );
buf_AQFP buf_splitterfromN146_n189_1_( clk_1 , splitterfromN146 , 0 , buf_splitterfromN146_n189_1 );
buf_AQFP buf_splitterfromN146_n189_2_( clk_3 , buf_splitterfromN146_n189_1 , 0 , buf_splitterfromN146_n189_2 );
buf_AQFP buf_splitterfromN146_n274_1_( clk_1 , splitterfromN146 , 0 , buf_splitterfromN146_n274_1 );
buf_AQFP buf_splitterfromN153_n148_1_( clk_8 , splitterfromN153 , 0 , buf_splitterfromN153_n148_1 );
buf_AQFP buf_splitterfromN153_n148_2_( clk_2 , buf_splitterfromN153_n148_1 , 0 , buf_splitterfromN153_n148_2 );
buf_AQFP buf_splitterfromN153_n290_1_( clk_8 , splitterfromN153 , 0 , buf_splitterfromN153_n290_1 );
buf_AQFP buf_splitterfromN153_n290_2_( clk_2 , buf_splitterfromN153_n290_1 , 0 , buf_splitterfromN153_n290_2 );
buf_AQFP buf_splitterN159ton117n330_n271_1_( clk_6 , splitterN159ton117n330 , 0 , buf_splitterN159ton117n330_n271_1 );
buf_AQFP buf_splitterN159ton117n330_n271_2_( clk_8 , buf_splitterN159ton117n330_n271_1 , 0 , buf_splitterN159ton117n330_n271_2 );
buf_AQFP buf_splitterN159ton117n330_n271_3_( clk_2 , buf_splitterN159ton117n330_n271_2 , 0 , buf_splitterN159ton117n330_n271_3 );
buf_AQFP buf_splitterN159ton117n330_n271_4_( clk_4 , buf_splitterN159ton117n330_n271_3 , 0 , buf_splitterN159ton117n330_n271_4 );
buf_AQFP buf_splitterN159ton117n330_n271_5_( clk_5 , buf_splitterN159ton117n330_n271_4 , 0 , buf_splitterN159ton117n330_n271_5 );
buf_AQFP buf_splitterN165ton129n346_n279_1_( clk_8 , splitterN165ton129n346 , 0 , buf_splitterN165ton129n346_n279_1 );
buf_AQFP buf_splitterN165ton129n346_n279_2_( clk_2 , buf_splitterN165ton129n346_n279_1 , 0 , buf_splitterN165ton129n346_n279_2 );
buf_AQFP buf_splitterN165ton129n346_n279_3_( clk_3 , buf_splitterN165ton129n346_n279_2 , 0 , buf_splitterN165ton129n346_n279_3 );
buf_AQFP buf_splitterN165ton129n346_n279_4_( clk_4 , buf_splitterN165ton129n346_n279_3 , 0 , buf_splitterN165ton129n346_n279_4 );
buf_AQFP buf_splitterN165ton129n346_n279_5_( clk_5 , buf_splitterN165ton129n346_n279_4 , 0 , buf_splitterN165ton129n346_n279_5 );
buf_AQFP buf_splitterN165ton280n346_n280_1_( clk_7 , splitterN165ton280n346 , 0 , buf_splitterN165ton280n346_n280_1 );
buf_AQFP buf_splitterN17ton146n68_n146_1_( clk_4 , splitterN17ton146n68 , 0 , buf_splitterN17ton146n68_n146_1 );
buf_AQFP buf_splitterN17ton146n68_n146_2_( clk_6 , buf_splitterN17ton146n68_n146_1 , 0 , buf_splitterN17ton146n68_n146_2 );
buf_AQFP buf_splitterN17ton146n68_n146_3_( clk_8 , buf_splitterN17ton146n68_n146_2 , 0 , buf_splitterN17ton146n68_n146_3 );
buf_AQFP buf_splitterN17ton159n68_n283_1_( clk_5 , splitterN17ton159n68 , 0 , buf_splitterN17ton159n68_n283_1 );
buf_AQFP buf_splitterN17ton159n68_n283_2_( clk_7 , buf_splitterN17ton159n68_n283_1 , 0 , buf_splitterN17ton159n68_n283_2 );
buf_AQFP buf_splitterN17ton159n68_n283_3_( clk_8 , buf_splitterN17ton159n68_n283_2 , 0 , buf_splitterN17ton159n68_n283_3 );
buf_AQFP buf_splitterN17ton159n68_n68_1_( clk_4 , splitterN17ton159n68 , 0 , buf_splitterN17ton159n68_n68_1 );
buf_AQFP buf_splitterN17ton159n68_n68_2_( clk_5 , buf_splitterN17ton159n68_n68_1 , 0 , buf_splitterN17ton159n68_n68_2 );
buf_AQFP buf_splitterN171ton132n361_n287_1_( clk_2 , splitterN171ton132n361 , 0 , buf_splitterN171ton132n361_n287_1 );
buf_AQFP buf_splitterN171ton132n361_n287_2_( clk_4 , buf_splitterN171ton132n361_n287_1 , 0 , buf_splitterN171ton132n361_n287_2 );
buf_AQFP buf_splitterN171ton132n361_n287_3_( clk_6 , buf_splitterN171ton132n361_n287_2 , 0 , buf_splitterN171ton132n361_n287_3 );
buf_AQFP buf_splitterN171ton288n361_n288_1_( clk_5 , splitterN171ton288n361 , 0 , buf_splitterN171ton288n361_n288_1 );
buf_AQFP buf_splitterN177ton117n315_n295_1_( clk_7 , splitterN177ton117n315 , 0 , buf_splitterN177ton117n315_n295_1 );
buf_AQFP buf_splitterN177ton117n315_n295_2_( clk_1 , buf_splitterN177ton117n315_n295_1 , 0 , buf_splitterN177ton117n315_n295_2 );
buf_AQFP buf_splitterN177ton117n315_n295_3_( clk_3 , buf_splitterN177ton117n315_n295_2 , 0 , buf_splitterN177ton117n315_n295_3 );
buf_AQFP buf_splitterN177ton117n315_n295_4_( clk_5 , buf_splitterN177ton117n315_n295_3 , 0 , buf_splitterN177ton117n315_n295_4 );
buf_AQFP buf_splitterN177ton296n315_n296_1_( clk_5 , splitterN177ton296n315 , 0 , buf_splitterN177ton296n315_n296_1 );
buf_AQFP buf_splitterN177ton296n315_n296_2_( clk_6 , buf_splitterN177ton296n315_n296_1 , 0 , buf_splitterN177ton296n315_n296_2 );
buf_AQFP buf_splitterN183ton132n221_n211_1_( clk_2 , splitterN183ton132n221 , 0 , buf_splitterN183ton132n221_n211_1 );
buf_AQFP buf_splitterN183ton132n221_n211_2_( clk_4 , buf_splitterN183ton132n221_n211_1 , 0 , buf_splitterN183ton132n221_n211_2 );
buf_AQFP buf_splitterN183ton132n221_n211_3_( clk_6 , buf_splitterN183ton132n221_n211_2 , 0 , buf_splitterN183ton132n221_n211_3 );
buf_AQFP buf_splitterN183ton212n221_n212_1_( clk_4 , splitterN183ton212n221 , 0 , buf_splitterN183ton212n221_n212_1 );
buf_AQFP buf_splitterN183ton212n221_n212_2_( clk_5 , buf_splitterN183ton212n221_n212_1 , 0 , buf_splitterN183ton212n221_n212_2 );
buf_AQFP buf_splitterN183ton212n221_n212_3_( clk_7 , buf_splitterN183ton212n221_n212_2 , 0 , buf_splitterN183ton212n221_n212_3 );
buf_AQFP buf_splitterN189ton123n236_n123_1_( clk_7 , splitterN189ton123n236 , 0 , buf_splitterN189ton123n236_n123_1 );
buf_AQFP buf_splitterN189ton123n236_n124_1_( clk_7 , splitterN189ton123n236 , 0 , buf_splitterN189ton123n236_n124_1 );
buf_AQFP buf_splitterN189ton123n236_n124_2_( clk_1 , buf_splitterN189ton123n236_n124_1 , 0 , buf_splitterN189ton123n236_n124_2 );
buf_AQFP buf_splitterN189ton123n236_n193_1_( clk_7 , splitterN189ton123n236 , 0 , buf_splitterN189ton123n236_n193_1 );
buf_AQFP buf_splitterN189ton123n236_n193_2_( clk_1 , buf_splitterN189ton123n236_n193_1 , 0 , buf_splitterN189ton123n236_n193_2 );
buf_AQFP buf_splitterN189ton123n236_n193_3_( clk_3 , buf_splitterN189ton123n236_n193_2 , 0 , buf_splitterN189ton123n236_n193_3 );
buf_AQFP buf_splitterN189ton123n236_n193_4_( clk_5 , buf_splitterN189ton123n236_n193_3 , 0 , buf_splitterN189ton123n236_n193_4 );
buf_AQFP buf_splitterN195ton123n253_n124_1_( clk_1 , splitterN195ton123n253 , 0 , buf_splitterN195ton123n253_n124_1 );
buf_AQFP buf_splitterN195ton123n253_n199_1_( clk_2 , splitterN195ton123n253 , 0 , buf_splitterN195ton123n253_n199_1 );
buf_AQFP buf_splitterN195ton123n253_n199_2_( clk_4 , buf_splitterN195ton123n253_n199_1 , 0 , buf_splitterN195ton123n253_n199_2 );
buf_AQFP buf_splitterN195ton123n253_n199_3_( clk_6 , buf_splitterN195ton123n253_n199_2 , 0 , buf_splitterN195ton123n253_n199_3 );
buf_AQFP buf_splitterN195ton200n253_n200_1_( clk_5 , splitterN195ton200n253 , 0 , buf_splitterN195ton200n253_n200_1 );
buf_AQFP buf_splitterN195ton200n253_n200_2_( clk_6 , buf_splitterN195ton200n253_n200_1 , 0 , buf_splitterN195ton200n253_n200_2 );
buf_AQFP buf_splitterN195ton200n253_n200_3_( clk_7 , buf_splitterN195ton200n253_n200_2 , 0 , buf_splitterN195ton200n253_n200_3 );
buf_AQFP buf_splitterN195ton200n253_n253_1_( clk_6 , splitterN195ton200n253 , 0 , buf_splitterN195ton200n253_n253_1 );
buf_AQFP buf_splitterN201ton129n180_n166_1_( clk_7 , splitterN201ton129n180 , 0 , buf_splitterN201ton129n180_n166_1 );
buf_AQFP buf_splitterN201ton129n180_n166_2_( clk_1 , buf_splitterN201ton129n180_n166_1 , 0 , buf_splitterN201ton129n180_n166_2 );
buf_AQFP buf_splitterN201ton129n180_n166_3_( clk_3 , buf_splitterN201ton129n180_n166_2 , 0 , buf_splitterN201ton129n180_n166_3 );
buf_AQFP buf_splitterN201ton129n180_n166_4_( clk_5 , buf_splitterN201ton129n180_n166_3 , 0 , buf_splitterN201ton129n180_n166_4 );
buf_AQFP buf_splitterN201ton167n180_n167_1_( clk_4 , splitterN201ton167n180 , 0 , buf_splitterN201ton167n180_n167_1 );
buf_AQFP buf_splitterN201ton167n180_n167_2_( clk_5 , buf_splitterN201ton167n180_n167_1 , 0 , buf_splitterN201ton167n180_n167_2 );
buf_AQFP buf_splitterN201ton167n180_n167_3_( clk_6 , buf_splitterN201ton167n180_n167_2 , 0 , buf_splitterN201ton167n180_n167_3 );
buf_AQFP buf_splitterN210ton182n360_n182_1_( clk_6 , splitterN210ton182n360 , 0 , buf_splitterN210ton182n360_n182_1 );
buf_AQFP buf_splitterN219ton171n355_n171_1_( clk_6 , splitterN219ton171n355 , 0 , buf_splitterN219ton171n355_n171_1 );
buf_AQFP buf_splitterN219ton171n355_n171_2_( clk_8 , buf_splitterN219ton171n355_n171_1 , 0 , buf_splitterN219ton171n355_n171_2 );
buf_AQFP buf_splitterN219ton171n355_n171_3_( clk_2 , buf_splitterN219ton171n355_n171_2 , 0 , buf_splitterN219ton171n355_n171_3 );
buf_AQFP buf_splitterN219ton171n355_n217_1_( clk_7 , splitterN219ton171n355 , 0 , buf_splitterN219ton171n355_n217_1 );
buf_AQFP buf_splitterN219ton171n355_n217_2_( clk_1 , buf_splitterN219ton171n355_n217_1 , 0 , buf_splitterN219ton171n355_n217_2 );
buf_AQFP buf_splitterN219ton171n355_n217_3_( clk_3 , buf_splitterN219ton171n355_n217_2 , 0 , buf_splitterN219ton171n355_n217_3 );
buf_AQFP buf_splitterN219ton171n355_n217_4_( clk_5 , buf_splitterN219ton171n355_n217_3 , 0 , buf_splitterN219ton171n355_n217_4 );
buf_AQFP buf_splitterN219ton171n355_n217_5_( clk_7 , buf_splitterN219ton171n355_n217_4 , 0 , buf_splitterN219ton171n355_n217_5 );
buf_AQFP buf_splitterN219ton171n355_n217_6_( clk_1 , buf_splitterN219ton171n355_n217_5 , 0 , buf_splitterN219ton171n355_n217_6 );
buf_AQFP buf_splitterN219ton171n355_n217_7_( clk_3 , buf_splitterN219ton171n355_n217_6 , 0 , buf_splitterN219ton171n355_n217_7 );
buf_AQFP buf_splitterN219ton232n308_n232_1_( clk_7 , splitterN219ton232n308 , 0 , buf_splitterN219ton232n308_n232_1 );
buf_AQFP buf_splitterN219ton232n308_n308_1_( clk_7 , splitterN219ton232n308 , 0 , buf_splitterN219ton232n308_n308_1 );
buf_AQFP buf_splitterN219ton232n308_n308_2_( clk_1 , buf_splitterN219ton232n308_n308_1 , 0 , buf_splitterN219ton232n308_n308_2 );
buf_AQFP buf_splitterN219ton232n308_n308_3_( clk_3 , buf_splitterN219ton232n308_n308_2 , 0 , buf_splitterN219ton232n308_n308_3 );
buf_AQFP buf_splitterN219ton232n308_n308_4_( clk_4 , buf_splitterN219ton232n308_n308_3 , 0 , buf_splitterN219ton232n308_n308_4 );
buf_AQFP buf_splitterN219ton311n355_n325_1_( clk_6 , splitterN219ton311n355 , 0 , buf_splitterN219ton311n355_n325_1 );
buf_AQFP buf_splitterN219ton311n355_n325_2_( clk_8 , buf_splitterN219ton311n355_n325_1 , 0 , buf_splitterN219ton311n355_n325_2 );
buf_AQFP buf_splitterN219ton311n355_n325_3_( clk_2 , buf_splitterN219ton311n355_n325_2 , 0 , buf_splitterN219ton311n355_n325_3 );
buf_AQFP buf_splitterN219ton311n355_n325_4_( clk_4 , buf_splitterN219ton311n355_n325_3 , 0 , buf_splitterN219ton311n355_n325_4 );
buf_AQFP buf_splitterN219ton311n355_n325_5_( clk_6 , buf_splitterN219ton311n355_n325_4 , 0 , buf_splitterN219ton311n355_n325_5 );
buf_AQFP buf_splitterN219ton311n355_n325_6_( clk_7 , buf_splitterN219ton311n355_n325_5 , 0 , buf_splitterN219ton311n355_n325_6 );
buf_AQFP buf_splitterN219ton311n355_n340_1_( clk_6 , splitterN219ton311n355 , 0 , buf_splitterN219ton311n355_n340_1 );
buf_AQFP buf_splitterN219ton311n355_n340_2_( clk_7 , buf_splitterN219ton311n355_n340_1 , 0 , buf_splitterN219ton311n355_n340_2 );
buf_AQFP buf_splitterN219ton311n355_n340_3_( clk_1 , buf_splitterN219ton311n355_n340_2 , 0 , buf_splitterN219ton311n355_n340_3 );
buf_AQFP buf_splitterN219ton311n355_n340_4_( clk_3 , buf_splitterN219ton311n355_n340_3 , 0 , buf_splitterN219ton311n355_n340_4 );
buf_AQFP buf_splitterN219ton311n355_n355_1_( clk_7 , splitterN219ton311n355 , 0 , buf_splitterN219ton311n355_n355_1 );
buf_AQFP buf_splitterN219ton311n355_n355_2_( clk_8 , buf_splitterN219ton311n355_n355_1 , 0 , buf_splitterN219ton311n355_n355_2 );
buf_AQFP buf_splitterN228ton173n357_n173_1_( clk_8 , splitterN228ton173n357 , 0 , buf_splitterN228ton173n357_n173_1 );
buf_AQFP buf_splitterN228ton173n357_n173_2_( clk_1 , buf_splitterN228ton173n357_n173_1 , 0 , buf_splitterN228ton173n357_n173_2 );
buf_AQFP buf_splitterN228ton173n357_n173_3_( clk_2 , buf_splitterN228ton173n357_n173_2 , 0 , buf_splitterN228ton173n357_n173_3 );
buf_AQFP buf_splitterN228ton173n357_n218_1_( clk_8 , splitterN228ton173n357 , 0 , buf_splitterN228ton173n357_n218_1 );
buf_AQFP buf_splitterN228ton173n357_n218_2_( clk_2 , buf_splitterN228ton173n357_n218_1 , 0 , buf_splitterN228ton173n357_n218_2 );
buf_AQFP buf_splitterN228ton309n357_n309_1_( clk_6 , splitterN228ton309n357 , 0 , buf_splitterN228ton309n357_n309_1 );
buf_AQFP buf_splitterN228ton309n357_n309_2_( clk_8 , buf_splitterN228ton309n357_n309_1 , 0 , buf_splitterN228ton309n357_n309_2 );
buf_AQFP buf_splitterN228ton309n357_n309_3_( clk_2 , buf_splitterN228ton309n357_n309_2 , 0 , buf_splitterN228ton309n357_n309_3 );
buf_AQFP buf_splitterN228ton309n357_n309_4_( clk_4 , buf_splitterN228ton309n357_n309_3 , 0 , buf_splitterN228ton309n357_n309_4 );
buf_AQFP buf_splitterN228ton309n357_n309_5_( clk_6 , buf_splitterN228ton309n357_n309_4 , 0 , buf_splitterN228ton309n357_n309_5 );
buf_AQFP buf_splitterN228ton309n357_n342_1_( clk_5 , splitterN228ton309n357 , 0 , buf_splitterN228ton309n357_n342_1 );
buf_AQFP buf_splitterN228ton309n357_n342_2_( clk_6 , buf_splitterN228ton309n357_n342_1 , 0 , buf_splitterN228ton309n357_n342_2 );
buf_AQFP buf_splitterN228ton309n357_n342_3_( clk_7 , buf_splitterN228ton309n357_n342_2 , 0 , buf_splitterN228ton309n357_n342_3 );
buf_AQFP buf_splitterN228ton309n357_n342_4_( clk_8 , buf_splitterN228ton309n357_n342_3 , 0 , buf_splitterN228ton309n357_n342_4 );
buf_AQFP buf_splitterN228ton309n357_n342_5_( clk_1 , buf_splitterN228ton309n357_n342_4 , 0 , buf_splitterN228ton309n357_n342_5 );
buf_AQFP buf_splitterN228ton309n357_n342_6_( clk_2 , buf_splitterN228ton309n357_n342_5 , 0 , buf_splitterN228ton309n357_n342_6 );
buf_AQFP buf_splitterN228ton309n357_n342_7_( clk_3 , buf_splitterN228ton309n357_n342_6 , 0 , buf_splitterN228ton309n357_n342_7 );
buf_AQFP buf_splitterN228ton309n357_n342_8_( clk_4 , buf_splitterN228ton309n357_n342_7 , 0 , buf_splitterN228ton309n357_n342_8 );
buf_AQFP buf_splitterN228ton309n357_n342_9_( clk_5 , buf_splitterN228ton309n357_n342_8 , 0 , buf_splitterN228ton309n357_n342_9 );
buf_AQFP buf_splitterN228ton309n357_n342_10_( clk_6 , buf_splitterN228ton309n357_n342_9 , 0 , buf_splitterN228ton309n357_n342_10 );
buf_AQFP buf_splitterN228ton309n357_n342_11_( clk_7 , buf_splitterN228ton309n357_n342_10 , 0 , buf_splitterN228ton309n357_n342_11 );
buf_AQFP buf_splitterN228ton309n357_n357_1_( clk_5 , splitterN228ton309n357 , 0 , buf_splitterN228ton309n357_n357_1 );
buf_AQFP buf_splitterN237ton174n358_n174_1_( clk_7 , splitterN237ton174n358 , 0 , buf_splitterN237ton174n358_n174_1 );
buf_AQFP buf_splitterN237ton174n358_n174_2_( clk_1 , buf_splitterN237ton174n358_n174_1 , 0 , buf_splitterN237ton174n358_n174_2 );
buf_AQFP buf_splitterN237ton174n358_n174_3_( clk_3 , buf_splitterN237ton174n358_n174_2 , 0 , buf_splitterN237ton174n358_n174_3 );
buf_AQFP buf_splitterN237ton174n358_n174_4_( clk_5 , buf_splitterN237ton174n358_n174_3 , 0 , buf_splitterN237ton174n358_n174_4 );
buf_AQFP buf_splitterN237ton174n358_n174_5_( clk_7 , buf_splitterN237ton174n358_n174_4 , 0 , buf_splitterN237ton174n358_n174_5 );
buf_AQFP buf_splitterN237ton174n358_n219_1_( clk_7 , splitterN237ton174n358 , 0 , buf_splitterN237ton174n358_n219_1 );
buf_AQFP buf_splitterN237ton174n358_n219_2_( clk_1 , buf_splitterN237ton174n358_n219_1 , 0 , buf_splitterN237ton174n358_n219_2 );
buf_AQFP buf_splitterN237ton174n358_n219_3_( clk_3 , buf_splitterN237ton174n358_n219_2 , 0 , buf_splitterN237ton174n358_n219_3 );
buf_AQFP buf_splitterN237ton174n358_n219_4_( clk_5 , buf_splitterN237ton174n358_n219_3 , 0 , buf_splitterN237ton174n358_n219_4 );
buf_AQFP buf_splitterN237ton174n358_n219_5_( clk_7 , buf_splitterN237ton174n358_n219_4 , 0 , buf_splitterN237ton174n358_n219_5 );
buf_AQFP buf_splitterN237ton174n358_n219_6_( clk_1 , buf_splitterN237ton174n358_n219_5 , 0 , buf_splitterN237ton174n358_n219_6 );
buf_AQFP buf_splitterN237ton313n358_n313_1_( clk_8 , splitterN237ton313n358 , 0 , buf_splitterN237ton313n358_n313_1 );
buf_AQFP buf_splitterN237ton313n358_n328_1_( clk_7 , splitterN237ton313n358 , 0 , buf_splitterN237ton313n358_n328_1 );
buf_AQFP buf_splitterN237ton313n358_n343_1_( clk_7 , splitterN237ton313n358 , 0 , buf_splitterN237ton313n358_n343_1 );
buf_AQFP buf_splitterN237ton313n358_n358_1_( clk_7 , splitterN237ton313n358 , 0 , buf_splitterN237ton313n358_n358_1 );
buf_AQFP buf_splitterN237ton313n358_n358_2_( clk_8 , buf_splitterN237ton313n358_n358_1 , 0 , buf_splitterN237ton313n358_n358_2 );
buf_AQFP buf_splitterN246ton175n359_n175_1_( clk_5 , splitterN246ton175n359 , 0 , buf_splitterN246ton175n359_n175_1 );
buf_AQFP buf_splitterN246ton175n359_n220_1_( clk_6 , splitterN246ton175n359 , 0 , buf_splitterN246ton175n359_n220_1 );
buf_AQFP buf_splitterN261ton169n201_n169_1_( clk_5 , splitterN261ton169n201 , 0 , buf_splitterN261ton169n201_n169_1 );
buf_AQFP buf_splitterN261ton169n201_n169_2_( clk_7 , buf_splitterN261ton169n201_n169_1 , 0 , buf_splitterN261ton169n201_n169_2 );
buf_AQFP buf_splitterN261ton169n201_n169_3_( clk_1 , buf_splitterN261ton169n201_n169_2 , 0 , buf_splitterN261ton169n201_n169_3 );
buf_AQFP buf_splitterN261ton169n201_n170_1_( clk_5 , splitterN261ton169n201 , 0 , buf_splitterN261ton169n201_n170_1 );
buf_AQFP buf_splitterN261ton169n201_n170_2_( clk_7 , buf_splitterN261ton169n201_n170_1 , 0 , buf_splitterN261ton169n201_n170_2 );
buf_AQFP buf_splitterN261ton169n201_n170_3_( clk_1 , buf_splitterN261ton169n201_n170_2 , 0 , buf_splitterN261ton169n201_n170_3 );
buf_AQFP buf_splitterN261ton169n201_n201_1_( clk_5 , splitterN261ton169n201 , 0 , buf_splitterN261ton169n201_n201_1 );
buf_AQFP buf_splitterN261ton169n201_n201_2_( clk_7 , buf_splitterN261ton169n201_n201_1 , 0 , buf_splitterN261ton169n201_n201_2 );
buf_AQFP buf_splitterN268ton152n331_n152_1_( clk_6 , splitterN268ton152n331 , 0 , buf_splitterN268ton152n331_n152_1 );
buf_AQFP buf_splitterN268ton152n331_n152_2_( clk_8 , buf_splitterN268ton152n331_n152_1 , 0 , buf_splitterN268ton152n331_n152_2 );
buf_AQFP buf_splitterN268ton152n331_n331_1_( clk_6 , splitterN268ton152n331 , 0 , buf_splitterN268ton152n331_n331_1 );
buf_AQFP buf_splitterN29ton61n84_n84_1_( clk_3 , splitterN29ton61n84 , 0 , buf_splitterN29ton61n84_n84_1 );
buf_AQFP buf_splitterN42ton153n77_n158_1_( clk_5 , splitterN42ton153n77 , 0 , buf_splitterN42ton153n77_n158_1 );
buf_AQFP buf_splitterN42ton176n77_n62_1_( clk_7 , splitterN42ton176n77 , 0 , buf_splitterN42ton176n77_n62_1 );
buf_AQFP buf_splitterN42ton176n77_n65_1_( clk_7 , splitterN42ton176n77 , 0 , buf_splitterN42ton176n77_n65_1 );
buf_AQFP buf_splitterN42ton176n77_n65_2_( clk_1 , buf_splitterN42ton176n77_n65_1 , 0 , buf_splitterN42ton176n77_n65_2 );
buf_AQFP buf_splitterN51ton159n81_n275_1_( clk_6 , splitterN51ton159n81 , 0 , buf_splitterN51ton159n81_n275_1 );
buf_AQFP buf_splitterN51ton159n81_n275_2_( clk_7 , buf_splitterN51ton159n81_n275_1 , 0 , buf_splitterN51ton159n81_n275_2 );
buf_AQFP buf_splitterN55ton151n82_n151_1_( clk_7 , splitterN55ton151n82 , 0 , buf_splitterN55ton151n82_n151_1 );
buf_AQFP buf_splitterN55ton151n82_n263_1_( clk_7 , splitterN55ton151n82 , 0 , buf_splitterN55ton151n82_n263_1 );
buf_AQFP buf_splitterN55ton151n82_n263_2_( clk_8 , buf_splitterN55ton151n82_n263_1 , 0 , buf_splitterN55ton151n82_n263_2 );
buf_AQFP buf_splitterfromN8_n267_1_( clk_3 , splitterfromN8 , 0 , buf_splitterfromN8_n267_1 );
buf_AQFP buf_splitterfromN8_n267_2_( clk_5 , buf_splitterfromN8_n267_1 , 0 , buf_splitterfromN8_n267_2 );
buf_AQFP buf_splitterfromN8_n267_3_( clk_7 , buf_splitterfromN8_n267_2 , 0 , buf_splitterfromN8_n267_3 );
buf_AQFP buf_splitterfromN8_n267_4_( clk_1 , buf_splitterfromN8_n267_3 , 0 , buf_splitterfromN8_n267_4 );
buf_AQFP buf_splitterN80ton149n76_n64_1_( clk_6 , splitterN80ton149n76 , 0 , buf_splitterN80ton149n76_n64_1 );
buf_AQFP buf_splitterN80ton149n76_n64_2_( clk_7 , buf_splitterN80ton149n76_n64_1 , 0 , buf_splitterN80ton149n76_n64_2 );
buf_AQFP buf_splitterN80ton149n76_n76_1_( clk_7 , splitterN80ton149n76 , 0 , buf_splitterN80ton149n76_n76_1 );
buf_AQFP buf_splitterN80ton149n76_n76_2_( clk_1 , buf_splitterN80ton149n76_n76_1 , 0 , buf_splitterN80ton149n76_n76_2 );
buf_AQFP buf_splitterN80ton149n76_n76_3_( clk_3 , buf_splitterN80ton149n76_n76_2 , 0 , buf_splitterN80ton149n76_n76_3 );
buf_AQFP buf_splitterN80ton149n76_n76_4_( clk_5 , buf_splitterN80ton149n76_n76_3 , 0 , buf_splitterN80ton149n76_n76_4 );
buf_AQFP buf_splitterN80ton149n76_n76_5_( clk_7 , buf_splitterN80ton149n76_n76_4 , 0 , buf_splitterN80ton149n76_n76_5 );
buf_AQFP buf_splitterN80ton149n76_n76_6_( clk_1 , buf_splitterN80ton149n76_n76_5 , 0 , buf_splitterN80ton149n76_n76_6 );
buf_AQFP buf_splitterN80ton149n76_n76_7_( clk_3 , buf_splitterN80ton149n76_n76_6 , 0 , buf_splitterN80ton149n76_n76_7 );
buf_AQFP buf_splitterN80ton149n76_n76_8_( clk_5 , buf_splitterN80ton149n76_n76_7 , 0 , buf_splitterN80ton149n76_n76_8 );
buf_AQFP buf_splitterN80ton149n76_n76_9_( clk_7 , buf_splitterN80ton149n76_n76_8 , 0 , buf_splitterN80ton149n76_n76_9 );
buf_AQFP buf_splitterN80ton149n76_n76_10_( clk_1 , buf_splitterN80ton149n76_n76_9 , 0 , buf_splitterN80ton149n76_n76_10 );
buf_AQFP buf_splitterN80ton149n76_n76_11_( clk_3 , buf_splitterN80ton149n76_n76_10 , 0 , buf_splitterN80ton149n76_n76_11 );
buf_AQFP buf_splitterN80ton149n76_n76_12_( clk_5 , buf_splitterN80ton149n76_n76_11 , 0 , buf_splitterN80ton149n76_n76_12 );
buf_AQFP buf_splitterN91ton262n94_n262_1_( clk_8 , splitterN91ton262n94 , 0 , buf_splitterN91ton262n94_n262_1 );
buf_AQFP buf_splitterN91ton262n94_n262_2_( clk_2 , buf_splitterN91ton262n94_n262_1 , 0 , buf_splitterN91ton262n94_n262_2 );
buf_AQFP buf_splitterN91ton262n94_n345_1_( clk_7 , splitterN91ton262n94 , 0 , buf_splitterN91ton262n94_n345_1 );
buf_AQFP buf_splitterN91ton262n94_n345_2_( clk_8 , buf_splitterN91ton262n94_n345_1 , 0 , buf_splitterN91ton262n94_n345_2 );
buf_AQFP buf_splitterN96ton273n91_n273_1_( clk_4 , splitterN96ton273n91 , 0 , buf_splitterN96ton273n91_n273_1 );
buf_AQFP buf_splitterN96ton273n91_n273_2_( clk_5 , buf_splitterN96ton273n91_n273_1 , 0 , buf_splitterN96ton273n91_n273_2 );
buf_AQFP buf_splitterN96ton273n91_n273_3_( clk_7 , buf_splitterN96ton273n91_n273_2 , 0 , buf_splitterN96ton273n91_n273_3 );
buf_AQFP buf_splitterN96ton273n91_n273_4_( clk_1 , buf_splitterN96ton273n91_n273_3 , 0 , buf_splitterN96ton273n91_n273_4 );
buf_AQFP buf_splitterN96ton273n91_n273_5_( clk_3 , buf_splitterN96ton273n91_n273_4 , 0 , buf_splitterN96ton273n91_n273_5 );
buf_AQFP buf_splitterN96ton273n91_n360_1_( clk_5 , splitterN96ton273n91 , 0 , buf_splitterN96ton273n91_n360_1 );
buf_AQFP buf_splitterN96ton273n91_n360_2_( clk_7 , buf_splitterN96ton273n91_n360_1 , 0 , buf_splitterN96ton273n91_n360_2 );
buf_AQFP buf_splitterfromn61_n62_1_( clk_7 , splitterfromn61 , 0 , buf_splitterfromn61_n62_1 );
buf_AQFP buf_splitterfromn63_n65_1_( clk_2 , splitterfromn63 , 0 , buf_splitterfromn63_n65_1 );
buf_AQFP buf_splittern65toN390n80_N390_1_( clk_4 , splittern65toN390n80 , 0 , buf_splittern65toN390n80_N390_1 );
buf_AQFP buf_splittern67ton160n83_n69_1_( clk_7 , splittern67ton160n83 , 0 , buf_splittern67ton160n83_n69_1 );
buf_AQFP buf_splittern67ton160n83_n69_2_( clk_1 , buf_splittern67ton160n83_n69_1 , 0 , buf_splittern67ton160n83_n69_2 );
buf_AQFP buf_splittern67ton160n83_n69_3_( clk_3 , buf_splittern67ton160n83_n69_2 , 0 , buf_splittern67ton160n83_n69_3 );
buf_AQFP buf_splittern67ton160n83_n69_4_( clk_5 , buf_splittern67ton160n83_n69_3 , 0 , buf_splittern67ton160n83_n69_4 );
buf_AQFP buf_splittern67ton160n83_n69_5_( clk_7 , buf_splittern67ton160n83_n69_4 , 0 , buf_splittern67ton160n83_n69_5 );
buf_AQFP buf_splittern67ton160n83_n69_6_( clk_1 , buf_splittern67ton160n83_n69_5 , 0 , buf_splittern67ton160n83_n69_6 );
buf_AQFP buf_splittern67ton160n83_n69_7_( clk_3 , buf_splittern67ton160n83_n69_6 , 0 , buf_splittern67ton160n83_n69_7 );
buf_AQFP buf_splittern67ton160n83_n69_8_( clk_5 , buf_splittern67ton160n83_n69_7 , 0 , buf_splittern67ton160n83_n69_8 );
buf_AQFP buf_splittern67ton160n83_n69_9_( clk_7 , buf_splittern67ton160n83_n69_8 , 0 , buf_splittern67ton160n83_n69_9 );
buf_AQFP buf_splittern67ton160n83_n69_10_( clk_1 , buf_splittern67ton160n83_n69_9 , 0 , buf_splittern67ton160n83_n69_10 );
buf_AQFP buf_splittern67ton160n83_n69_11_( clk_3 , buf_splittern67ton160n83_n69_10 , 0 , buf_splittern67ton160n83_n69_11 );
buf_AQFP buf_splittern67ton160n83_n83_1_( clk_7 , splittern67ton160n83 , 0 , buf_splittern67ton160n83_n83_1 );
buf_AQFP buf_splitterfromn68_n69_1_( clk_3 , splitterfromn68 , 0 , buf_splitterfromn68_n69_1 );
buf_AQFP buf_splitterfromn68_n69_2_( clk_4 , buf_splitterfromn68_n69_1 , 0 , buf_splitterfromn68_n69_2 );
buf_AQFP buf_splitterfromn68_n69_3_( clk_5 , buf_splitterfromn68_n69_2 , 0 , buf_splitterfromn68_n69_3 );
buf_AQFP buf_splitterfromn68_n69_4_( clk_7 , buf_splitterfromn68_n69_3 , 0 , buf_splitterfromn68_n69_4 );
buf_AQFP buf_splitterfromn68_n69_5_( clk_1 , buf_splitterfromn68_n69_4 , 0 , buf_splitterfromn68_n69_5 );
buf_AQFP buf_splitterfromn68_n69_6_( clk_3 , buf_splitterfromn68_n69_5 , 0 , buf_splitterfromn68_n69_6 );
buf_AQFP buf_splitterfromn68_n71_1_( clk_3 , splitterfromn68 , 0 , buf_splitterfromn68_n71_1 );
buf_AQFP buf_splitterfromn68_n71_2_( clk_5 , buf_splitterfromn68_n71_1 , 0 , buf_splitterfromn68_n71_2 );
buf_AQFP buf_splitterfromn68_n71_3_( clk_7 , buf_splitterfromn68_n71_2 , 0 , buf_splitterfromn68_n71_3 );
buf_AQFP buf_splitterfromn68_n71_4_( clk_1 , buf_splitterfromn68_n71_3 , 0 , buf_splitterfromn68_n71_4 );
buf_AQFP buf_splitterfromn70_n71_1_( clk_5 , splitterfromn70 , 0 , buf_splitterfromn70_n71_1 );
buf_AQFP buf_splitterfromn70_n71_2_( clk_6 , buf_splitterfromn70_n71_1 , 0 , buf_splitterfromn70_n71_2 );
buf_AQFP buf_splitterfromn70_n71_3_( clk_8 , buf_splitterfromn70_n71_2 , 0 , buf_splitterfromn70_n71_3 );
buf_AQFP buf_splitterfromn70_n71_4_( clk_2 , buf_splitterfromn70_n71_3 , 0 , buf_splitterfromn70_n71_4 );
buf_AQFP buf_splitterfromn70_n71_5_( clk_4 , buf_splitterfromn70_n71_4 , 0 , buf_splitterfromn70_n71_5 );
buf_AQFP buf_splitterfromn70_n71_6_( clk_6 , buf_splitterfromn70_n71_5 , 0 , buf_splitterfromn70_n71_6 );
buf_AQFP buf_splitterfromn70_n71_7_( clk_8 , buf_splitterfromn70_n71_6 , 0 , buf_splitterfromn70_n71_7 );
buf_AQFP buf_splitterfromn70_n71_8_( clk_2 , buf_splitterfromn70_n71_7 , 0 , buf_splitterfromn70_n71_8 );
buf_AQFP buf_splitterfromn70_n71_9_( clk_4 , buf_splitterfromn70_n71_8 , 0 , buf_splitterfromn70_n71_9 );
buf_AQFP buf_splitterfromn70_n71_10_( clk_6 , buf_splitterfromn70_n71_9 , 0 , buf_splitterfromn70_n71_10 );
buf_AQFP buf_splitterfromn70_n71_11_( clk_8 , buf_splitterfromn70_n71_10 , 0 , buf_splitterfromn70_n71_11 );
buf_AQFP buf_splitterfromn70_n71_12_( clk_2 , buf_splitterfromn70_n71_11 , 0 , buf_splitterfromn70_n71_12 );
buf_AQFP buf_splitterfromn71_n72_1_( clk_1 , splitterfromn71 , 0 , buf_splitterfromn71_n72_1 );
buf_AQFP buf_splitterfromn71_n80_1_( clk_1 , splitterfromn71 , 0 , buf_splitterfromn71_n80_1 );
buf_AQFP buf_splitterfromn75_n76_1_( clk_6 , splitterfromn75 , 0 , buf_splitterfromn75_n76_1 );
buf_AQFP buf_splitterfromn75_n76_2_( clk_8 , buf_splitterfromn75_n76_1 , 0 , buf_splitterfromn75_n76_2 );
buf_AQFP buf_splitterfromn75_n76_3_( clk_2 , buf_splitterfromn75_n76_2 , 0 , buf_splitterfromn75_n76_3 );
buf_AQFP buf_splitterfromn75_n76_4_( clk_4 , buf_splitterfromn75_n76_3 , 0 , buf_splitterfromn75_n76_4 );
buf_AQFP buf_splitterfromn75_n76_5_( clk_6 , buf_splitterfromn75_n76_4 , 0 , buf_splitterfromn75_n76_5 );
buf_AQFP buf_splitterfromn75_n76_6_( clk_8 , buf_splitterfromn75_n76_5 , 0 , buf_splitterfromn75_n76_6 );
buf_AQFP buf_splitterfromn75_n76_7_( clk_2 , buf_splitterfromn75_n76_6 , 0 , buf_splitterfromn75_n76_7 );
buf_AQFP buf_splitterfromn75_n76_8_( clk_4 , buf_splitterfromn75_n76_7 , 0 , buf_splitterfromn75_n76_8 );
buf_AQFP buf_splitterfromn75_n76_9_( clk_6 , buf_splitterfromn75_n76_8 , 0 , buf_splitterfromn75_n76_9 );
buf_AQFP buf_splitterfromn75_n76_10_( clk_8 , buf_splitterfromn75_n76_9 , 0 , buf_splitterfromn75_n76_10 );
buf_AQFP buf_splitterfromn75_n76_11_( clk_2 , buf_splitterfromn75_n76_10 , 0 , buf_splitterfromn75_n76_11 );
buf_AQFP buf_splitterfromn75_n76_12_( clk_4 , buf_splitterfromn75_n76_11 , 0 , buf_splitterfromn75_n76_12 );
buf_AQFP buf_splitterfromn75_n76_13_( clk_6 , buf_splitterfromn75_n76_12 , 0 , buf_splitterfromn75_n76_13 );
buf_AQFP buf_splitterfromn78_n79_1_( clk_6 , splitterfromn78 , 0 , buf_splitterfromn78_n79_1 );
buf_AQFP buf_splitterfromn78_n79_2_( clk_8 , buf_splitterfromn78_n79_1 , 0 , buf_splitterfromn78_n79_2 );
buf_AQFP buf_splitterfromn78_n89_1_( clk_6 , splitterfromn78 , 0 , buf_splitterfromn78_n89_1 );
buf_AQFP buf_splittern81toN447n156_N447_1_( clk_8 , splittern81toN447n156 , 0 , buf_splittern81toN447n156_N447_1 );
buf_AQFP buf_splittern81toN447n156_N447_2_( clk_2 , buf_splittern81toN447n156_N447_1 , 0 , buf_splittern81toN447n156_N447_2 );
buf_AQFP buf_splittern81toN447n156_N447_3_( clk_4 , buf_splittern81toN447n156_N447_2 , 0 , buf_splittern81toN447n156_N447_3 );
buf_AQFP buf_splittern81toN447n156_N447_4_( clk_6 , buf_splittern81toN447n156_N447_3 , 0 , buf_splittern81toN447n156_N447_4 );
buf_AQFP buf_splittern81toN447n156_N447_5_( clk_8 , buf_splittern81toN447n156_N447_4 , 0 , buf_splittern81toN447n156_N447_5 );
buf_AQFP buf_splittern81toN447n156_N447_6_( clk_2 , buf_splittern81toN447n156_N447_5 , 0 , buf_splittern81toN447n156_N447_6 );
buf_AQFP buf_splittern81toN447n156_N447_7_( clk_4 , buf_splittern81toN447n156_N447_6 , 0 , buf_splittern81toN447n156_N447_7 );
buf_AQFP buf_splittern81toN447n156_N447_8_( clk_6 , buf_splittern81toN447n156_N447_7 , 0 , buf_splittern81toN447n156_N447_8 );
buf_AQFP buf_splittern81toN447n156_N447_9_( clk_8 , buf_splittern81toN447n156_N447_8 , 0 , buf_splittern81toN447n156_N447_9 );
buf_AQFP buf_splittern81toN447n156_N447_10_( clk_2 , buf_splittern81toN447n156_N447_9 , 0 , buf_splittern81toN447n156_N447_10 );
buf_AQFP buf_splittern81toN447n156_N447_11_( clk_4 , buf_splittern81toN447n156_N447_10 , 0 , buf_splittern81toN447n156_N447_11 );
buf_AQFP buf_splittern81toN447n156_N447_12_( clk_6 , buf_splittern81toN447n156_N447_11 , 0 , buf_splittern81toN447n156_N447_12 );
buf_AQFP buf_splittern81toN447n156_N447_13_( clk_8 , buf_splittern81toN447n156_N447_12 , 0 , buf_splittern81toN447n156_N447_13 );
buf_AQFP buf_splittern81toN447n156_N447_14_( clk_2 , buf_splittern81toN447n156_N447_13 , 0 , buf_splittern81toN447n156_N447_14 );
buf_AQFP buf_splittern81toN447n156_N447_15_( clk_4 , buf_splittern81toN447n156_N447_14 , 0 , buf_splittern81toN447n156_N447_15 );
buf_AQFP buf_splittern81toN447n156_N447_16_( clk_6 , buf_splittern81toN447n156_N447_15 , 0 , buf_splittern81toN447n156_N447_16 );
buf_AQFP buf_splittern81toN447n156_N447_17_( clk_7 , buf_splittern81toN447n156_N447_16 , 0 , buf_splittern81toN447n156_N447_17 );
buf_AQFP buf_splittern81toN447n156_N447_18_( clk_1 , buf_splittern81toN447n156_N447_17 , 0 , buf_splittern81toN447n156_N447_18 );
buf_AQFP buf_splittern81toN447n156_N447_19_( clk_3 , buf_splittern81toN447n156_N447_18 , 0 , buf_splittern81toN447n156_N447_19 );
buf_AQFP buf_splittern83ton179n88_n85_1_( clk_3 , splittern83ton179n88 , 0 , buf_splittern83ton179n88_n85_1 );
buf_AQFP buf_splittern83ton179n88_n85_2_( clk_5 , buf_splittern83ton179n88_n85_1 , 0 , buf_splittern83ton179n88_n85_2 );
buf_AQFP buf_splittern83ton179n88_n85_3_( clk_7 , buf_splittern83ton179n88_n85_2 , 0 , buf_splittern83ton179n88_n85_3 );
buf_AQFP buf_splittern83ton179n88_n85_4_( clk_1 , buf_splittern83ton179n88_n85_3 , 0 , buf_splittern83ton179n88_n85_4 );
buf_AQFP buf_splittern83ton179n88_n85_5_( clk_3 , buf_splittern83ton179n88_n85_4 , 0 , buf_splittern83ton179n88_n85_5 );
buf_AQFP buf_splittern83ton179n88_n85_6_( clk_4 , buf_splittern83ton179n88_n85_5 , 0 , buf_splittern83ton179n88_n85_6 );
buf_AQFP buf_splittern83ton179n88_n85_7_( clk_5 , buf_splittern83ton179n88_n85_6 , 0 , buf_splittern83ton179n88_n85_7 );
buf_AQFP buf_splittern83ton179n88_n85_8_( clk_7 , buf_splittern83ton179n88_n85_7 , 0 , buf_splittern83ton179n88_n85_8 );
buf_AQFP buf_splittern83ton179n88_n85_9_( clk_8 , buf_splittern83ton179n88_n85_8 , 0 , buf_splittern83ton179n88_n85_9 );
buf_AQFP buf_splittern83ton179n88_n85_10_( clk_2 , buf_splittern83ton179n88_n85_9 , 0 , buf_splittern83ton179n88_n85_10 );
buf_AQFP buf_splittern83ton179n88_n85_11_( clk_4 , buf_splittern83ton179n88_n85_10 , 0 , buf_splittern83ton179n88_n85_11 );
buf_AQFP buf_splittern83ton179n88_n85_12_( clk_6 , buf_splittern83ton179n88_n85_11 , 0 , buf_splittern83ton179n88_n85_12 );
buf_AQFP buf_splittern83ton179n88_n85_13_( clk_7 , buf_splittern83ton179n88_n85_12 , 0 , buf_splittern83ton179n88_n85_13 );
buf_AQFP buf_splittern83ton179n88_n85_14_( clk_8 , buf_splittern83ton179n88_n85_13 , 0 , buf_splittern83ton179n88_n85_14 );
buf_AQFP buf_splittern83ton179n88_n85_15_( clk_2 , buf_splittern83ton179n88_n85_14 , 0 , buf_splittern83ton179n88_n85_15 );
buf_AQFP buf_splittern83ton179n88_n85_16_( clk_4 , buf_splittern83ton179n88_n85_15 , 0 , buf_splittern83ton179n88_n85_16 );
buf_AQFP buf_splitterfromn95_n114_1_( clk_5 , splitterfromn95 , 0 , buf_splitterfromn95_n114_1 );
buf_AQFP buf_splitterfromn95_n114_2_( clk_7 , buf_splitterfromn95_n114_1 , 0 , buf_splitterfromn95_n114_2 );
buf_AQFP buf_splitterfromn95_n114_3_( clk_1 , buf_splitterfromn95_n114_2 , 0 , buf_splitterfromn95_n114_3 );
buf_AQFP buf_splitterfromn95_n114_4_( clk_3 , buf_splitterfromn95_n114_3 , 0 , buf_splitterfromn95_n114_4 );
buf_AQFP buf_splitterfromn95_n114_5_( clk_5 , buf_splitterfromn95_n114_4 , 0 , buf_splitterfromn95_n114_5 );
buf_AQFP buf_splitterfromn95_n114_6_( clk_7 , buf_splitterfromn95_n114_5 , 0 , buf_splitterfromn95_n114_6 );
buf_AQFP buf_splitterfromn95_n114_7_( clk_8 , buf_splitterfromn95_n114_6 , 0 , buf_splitterfromn95_n114_7 );
buf_AQFP buf_splitterfromn95_n114_8_( clk_1 , buf_splitterfromn95_n114_7 , 0 , buf_splitterfromn95_n114_8 );
buf_AQFP buf_splitterfromn95_n114_9_( clk_2 , buf_splitterfromn95_n114_8 , 0 , buf_splitterfromn95_n114_9 );
buf_AQFP buf_splitterfromn95_n114_10_( clk_3 , buf_splitterfromn95_n114_9 , 0 , buf_splitterfromn95_n114_10 );
buf_AQFP buf_splitterfromn95_n114_11_( clk_5 , buf_splitterfromn95_n114_10 , 0 , buf_splitterfromn95_n114_11 );
buf_AQFP buf_splitterfromn95_n114_12_( clk_7 , buf_splitterfromn95_n114_11 , 0 , buf_splitterfromn95_n114_12 );
buf_AQFP buf_splitterfromn95_n115_1_( clk_5 , splitterfromn95 , 0 , buf_splitterfromn95_n115_1 );
buf_AQFP buf_splitterfromn95_n115_2_( clk_7 , buf_splitterfromn95_n115_1 , 0 , buf_splitterfromn95_n115_2 );
buf_AQFP buf_splitterfromn95_n115_3_( clk_8 , buf_splitterfromn95_n115_2 , 0 , buf_splitterfromn95_n115_3 );
buf_AQFP buf_splitterfromn95_n115_4_( clk_2 , buf_splitterfromn95_n115_3 , 0 , buf_splitterfromn95_n115_4 );
buf_AQFP buf_splitterfromn95_n115_5_( clk_3 , buf_splitterfromn95_n115_4 , 0 , buf_splitterfromn95_n115_5 );
buf_AQFP buf_splitterfromn95_n115_6_( clk_4 , buf_splitterfromn95_n115_5 , 0 , buf_splitterfromn95_n115_6 );
buf_AQFP buf_splitterfromn95_n115_7_( clk_5 , buf_splitterfromn95_n115_6 , 0 , buf_splitterfromn95_n115_7 );
buf_AQFP buf_splitterfromn95_n115_8_( clk_6 , buf_splitterfromn95_n115_7 , 0 , buf_splitterfromn95_n115_8 );
buf_AQFP buf_splitterfromn104_n109_1_( clk_2 , splitterfromn104 , 0 , buf_splitterfromn104_n109_1 );
buf_AQFP buf_splitterfromn113_n114_1_( clk_7 , splitterfromn113 , 0 , buf_splitterfromn113_n114_1 );
buf_AQFP buf_splitterfromn113_n114_2_( clk_8 , buf_splitterfromn113_n114_1 , 0 , buf_splitterfromn113_n114_2 );
buf_AQFP buf_splitterfromn113_n114_3_( clk_1 , buf_splitterfromn113_n114_2 , 0 , buf_splitterfromn113_n114_3 );
buf_AQFP buf_splitterfromn113_n114_4_( clk_3 , buf_splitterfromn113_n114_3 , 0 , buf_splitterfromn113_n114_4 );
buf_AQFP buf_splitterfromn113_n114_5_( clk_5 , buf_splitterfromn113_n114_4 , 0 , buf_splitterfromn113_n114_5 );
buf_AQFP buf_splitterfromn113_n114_6_( clk_7 , buf_splitterfromn113_n114_5 , 0 , buf_splitterfromn113_n114_6 );
buf_AQFP buf_splitterfromn113_n114_7_( clk_1 , buf_splitterfromn113_n114_6 , 0 , buf_splitterfromn113_n114_7 );
buf_AQFP buf_splitterfromn113_n114_8_( clk_3 , buf_splitterfromn113_n114_7 , 0 , buf_splitterfromn113_n114_8 );
buf_AQFP buf_splitterfromn113_n114_9_( clk_4 , buf_splitterfromn113_n114_8 , 0 , buf_splitterfromn113_n114_9 );
buf_AQFP buf_splitterfromn113_n114_10_( clk_5 , buf_splitterfromn113_n114_9 , 0 , buf_splitterfromn113_n114_10 );
buf_AQFP buf_splitterfromn113_n114_11_( clk_6 , buf_splitterfromn113_n114_10 , 0 , buf_splitterfromn113_n114_11 );
buf_AQFP buf_splitterfromn113_n114_12_( clk_7 , buf_splitterfromn113_n114_11 , 0 , buf_splitterfromn113_n114_12 );
buf_AQFP buf_splitterfromn113_n114_13_( clk_8 , buf_splitterfromn113_n114_12 , 0 , buf_splitterfromn113_n114_13 );
buf_AQFP buf_splitterfromn113_n115_1_( clk_8 , splitterfromn113 , 0 , buf_splitterfromn113_n115_1 );
buf_AQFP buf_splitterfromn113_n115_2_( clk_2 , buf_splitterfromn113_n115_1 , 0 , buf_splitterfromn113_n115_2 );
buf_AQFP buf_splitterfromn113_n115_3_( clk_3 , buf_splitterfromn113_n115_2 , 0 , buf_splitterfromn113_n115_3 );
buf_AQFP buf_splitterfromn113_n115_4_( clk_4 , buf_splitterfromn113_n115_3 , 0 , buf_splitterfromn113_n115_4 );
buf_AQFP buf_splitterfromn113_n115_5_( clk_6 , buf_splitterfromn113_n115_4 , 0 , buf_splitterfromn113_n115_5 );
buf_AQFP buf_splitterfromn122_n141_1_( clk_8 , splitterfromn122 , 0 , buf_splitterfromn122_n141_1 );
buf_AQFP buf_splitterfromn122_n142_1_( clk_7 , splitterfromn122 , 0 , buf_splitterfromn122_n142_1 );
buf_AQFP buf_splitterfromn122_n142_2_( clk_8 , buf_splitterfromn122_n142_1 , 0 , buf_splitterfromn122_n142_2 );
buf_AQFP buf_splitterfromn122_n142_3_( clk_1 , buf_splitterfromn122_n142_2 , 0 , buf_splitterfromn122_n142_3 );
buf_AQFP buf_splitterfromn131_n136_1_( clk_4 , splitterfromn131 , 0 , buf_splitterfromn131_n136_1 );
buf_AQFP buf_splitterfromn134_n136_1_( clk_4 , splitterfromn134 , 0 , buf_splitterfromn134_n136_1 );
buf_AQFP buf_splitterfromn144_n145_1_( clk_6 , splitterfromn144 , 0 , buf_splitterfromn144_n145_1 );
buf_AQFP buf_splitterfromn144_n156_1_( clk_5 , splitterfromn144 , 0 , buf_splitterfromn144_n156_1 );
buf_AQFP buf_splittern152ton164n210_n210_1_( clk_4 , splittern152ton164n210 , 0 , buf_splittern152ton164n210_n210_1 );
buf_AQFP buf_splittern152ton164n210_n210_2_( clk_5 , buf_splittern152ton164n210_n210_1 , 0 , buf_splittern152ton164n210_n210_2 );
buf_AQFP buf_splittern193ton206n234_n206_1_( clk_1 , splittern193ton206n234 , 0 , buf_splittern193ton206n234_n206_1 );
buf_AQFP buf_splittern193ton206n234_n206_2_( clk_3 , buf_splittern193ton206n234_n206_1 , 0 , buf_splittern193ton206n234_n206_2 );
buf_AQFP buf_splittern193ton206n234_n206_3_( clk_5 , buf_splittern193ton206n234_n206_2 , 0 , buf_splittern193ton206n234_n206_3 );
buf_AQFP buf_splittern193ton206n234_n206_4_( clk_6 , buf_splittern193ton206n234_n206_3 , 0 , buf_splittern193ton206n234_n206_4 );
buf_AQFP buf_splitterfromn194_n205_1_( clk_2 , splitterfromn194 , 0 , buf_splitterfromn194_n205_1 );
buf_AQFP buf_splitterfromn194_n205_2_( clk_4 , buf_splitterfromn194_n205_1 , 0 , buf_splitterfromn194_n205_2 );
buf_AQFP buf_splitterfromn194_n205_3_( clk_5 , buf_splitterfromn194_n205_2 , 0 , buf_splitterfromn194_n205_3 );
buf_AQFP buf_splittern199ton204n251_n204_1_( clk_3 , splittern199ton204n251 , 0 , buf_splittern199ton204n251_n204_1 );
buf_AQFP buf_splitterfromn200_n203_1_( clk_2 , splitterfromn200 , 0 , buf_splitterfromn200_n203_1 );
buf_AQFP buf_splittern211ton213n298_n298_1_( clk_3 , splittern211ton213n298 , 0 , buf_splittern211ton213n298_n298_1 );
buf_AQFP buf_splittern211ton213n298_n298_2_( clk_5 , buf_splittern211ton213n298_n298_1 , 0 , buf_splittern211ton213n298_n298_2 );
buf_AQFP buf_splittern211ton213n298_n298_3_( clk_7 , buf_splittern211ton213n298_n298_2 , 0 , buf_splittern211ton213n298_n298_3 );
buf_AQFP buf_splittern211ton213n298_n298_4_( clk_1 , buf_splittern211ton213n298_n298_3 , 0 , buf_splittern211ton213n298_n298_4 );
buf_AQFP buf_splitterfromn212_n297_1_( clk_3 , splitterfromn212 , 0 , buf_splitterfromn212_n297_1 );
buf_AQFP buf_splitterfromn212_n297_2_( clk_5 , buf_splitterfromn212_n297_1 , 0 , buf_splitterfromn212_n297_2 );
buf_AQFP buf_splitterfromn212_n297_3_( clk_6 , buf_splitterfromn212_n297_2 , 0 , buf_splitterfromn212_n297_3 );
buf_AQFP buf_splitterfromn212_n297_4_( clk_7 , buf_splitterfromn212_n297_3 , 0 , buf_splitterfromn212_n297_4 );
buf_AQFP buf_splitterfromn212_n297_5_( clk_8 , buf_splitterfromn212_n297_4 , 0 , buf_splitterfromn212_n297_5 );
buf_AQFP buf_splitterfromn212_n297_6_( clk_1 , buf_splitterfromn212_n297_5 , 0 , buf_splitterfromn212_n297_6 );
buf_AQFP buf_splittern213ton214n218_n214_1_( clk_5 , splittern213ton214n218 , 0 , buf_splittern213ton214n218_n214_1 );
buf_AQFP buf_splittern213ton214n218_n214_2_( clk_6 , buf_splittern213ton214n218_n214_1 , 0 , buf_splittern213ton214n218_n214_2 );
buf_AQFP buf_splittern213ton214n218_n214_3_( clk_8 , buf_splittern213ton214n218_n214_2 , 0 , buf_splittern213ton214n218_n214_3 );
buf_AQFP buf_splittern213ton214n218_n215_1_( clk_5 , splittern213ton214n218 , 0 , buf_splittern213ton214n218_n215_1 );
buf_AQFP buf_splittern213ton214n218_n215_2_( clk_6 , buf_splittern213ton214n218_n215_1 , 0 , buf_splittern213ton214n218_n215_2 );
buf_AQFP buf_splittern213ton214n218_n215_3_( clk_8 , buf_splittern213ton214n218_n215_2 , 0 , buf_splittern213ton214n218_n215_3 );
buf_AQFP buf_splittern228ton229n233_n229_1_( clk_4 , splittern228ton229n233 , 0 , buf_splittern228ton229n233_n229_1 );
buf_AQFP buf_splittern228ton229n233_n229_2_( clk_6 , buf_splittern228ton229n233_n229_1 , 0 , buf_splittern228ton229n233_n229_2 );
buf_AQFP buf_splittern228ton229n233_n230_1_( clk_4 , splittern228ton229n233 , 0 , buf_splittern228ton229n233_n230_1 );
buf_AQFP buf_splittern228ton229n233_n230_2_( clk_6 , buf_splittern228ton229n233_n230_1 , 0 , buf_splittern228ton229n233_n230_2 );
buf_AQFP buf_splittern271ton306n328_n306_1_( clk_1 , splittern271ton306n328 , 0 , buf_splittern271ton306n328_n306_1 );
buf_AQFP buf_splittern271ton306n328_n306_2_( clk_3 , buf_splittern271ton306n328_n306_1 , 0 , buf_splittern271ton306n328_n306_2 );
buf_AQFP buf_splittern271ton306n328_n306_3_( clk_5 , buf_splittern271ton306n328_n306_2 , 0 , buf_splittern271ton306n328_n306_3 );
buf_AQFP buf_splittern271ton306n328_n306_4_( clk_7 , buf_splittern271ton306n328_n306_3 , 0 , buf_splittern271ton306n328_n306_4 );
buf_AQFP buf_splittern271ton306n328_n306_5_( clk_1 , buf_splittern271ton306n328_n306_4 , 0 , buf_splittern271ton306n328_n306_5 );
buf_AQFP buf_splittern271ton306n328_n306_6_( clk_2 , buf_splittern271ton306n328_n306_5 , 0 , buf_splittern271ton306n328_n306_6 );
buf_AQFP buf_splittern271ton306n328_n306_7_( clk_4 , buf_splittern271ton306n328_n306_6 , 0 , buf_splittern271ton306n328_n306_7 );
buf_AQFP buf_splittern271ton306n328_n306_8_( clk_6 , buf_splittern271ton306n328_n306_7 , 0 , buf_splittern271ton306n328_n306_8 );
buf_AQFP buf_splittern271ton306n328_n306_9_( clk_8 , buf_splittern271ton306n328_n306_8 , 0 , buf_splittern271ton306n328_n306_9 );
buf_AQFP buf_splittern271ton306n328_n306_10_( clk_2 , buf_splittern271ton306n328_n306_9 , 0 , buf_splittern271ton306n328_n306_10 );
buf_AQFP buf_splittern271ton306n328_n306_11_( clk_4 , buf_splittern271ton306n328_n306_10 , 0 , buf_splittern271ton306n328_n306_11 );
buf_AQFP buf_splittern271ton306n328_n306_12_( clk_6 , buf_splittern271ton306n328_n306_11 , 0 , buf_splittern271ton306n328_n306_12 );
buf_AQFP buf_splitterfromn272_n305_1_( clk_3 , splitterfromn272 , 0 , buf_splitterfromn272_n305_1 );
buf_AQFP buf_splitterfromn272_n305_2_( clk_5 , buf_splitterfromn272_n305_1 , 0 , buf_splitterfromn272_n305_2 );
buf_AQFP buf_splitterfromn272_n305_3_( clk_7 , buf_splitterfromn272_n305_2 , 0 , buf_splitterfromn272_n305_3 );
buf_AQFP buf_splitterfromn272_n305_4_( clk_1 , buf_splitterfromn272_n305_3 , 0 , buf_splitterfromn272_n305_4 );
buf_AQFP buf_splitterfromn272_n305_5_( clk_3 , buf_splitterfromn272_n305_4 , 0 , buf_splitterfromn272_n305_5 );
buf_AQFP buf_splitterfromn272_n305_6_( clk_5 , buf_splitterfromn272_n305_5 , 0 , buf_splitterfromn272_n305_6 );
buf_AQFP buf_splitterfromn272_n305_7_( clk_7 , buf_splitterfromn272_n305_6 , 0 , buf_splitterfromn272_n305_7 );
buf_AQFP buf_splitterfromn272_n305_8_( clk_1 , buf_splitterfromn272_n305_7 , 0 , buf_splitterfromn272_n305_8 );
buf_AQFP buf_splitterfromn272_n305_9_( clk_2 , buf_splitterfromn272_n305_8 , 0 , buf_splitterfromn272_n305_9 );
buf_AQFP buf_splitterfromn272_n305_10_( clk_4 , buf_splitterfromn272_n305_9 , 0 , buf_splitterfromn272_n305_10 );
buf_AQFP buf_splittern279ton304n343_n304_1_( clk_2 , splittern279ton304n343 , 0 , buf_splittern279ton304n343_n304_1 );
buf_AQFP buf_splittern279ton304n343_n304_2_( clk_4 , buf_splittern279ton304n343_n304_1 , 0 , buf_splittern279ton304n343_n304_2 );
buf_AQFP buf_splittern279ton304n343_n304_3_( clk_6 , buf_splittern279ton304n343_n304_2 , 0 , buf_splittern279ton304n343_n304_3 );
buf_AQFP buf_splittern279ton304n343_n304_4_( clk_8 , buf_splittern279ton304n343_n304_3 , 0 , buf_splittern279ton304n343_n304_4 );
buf_AQFP buf_splittern279ton304n343_n304_5_( clk_2 , buf_splittern279ton304n343_n304_4 , 0 , buf_splittern279ton304n343_n304_5 );
buf_AQFP buf_splittern279ton304n343_n304_6_( clk_4 , buf_splittern279ton304n343_n304_5 , 0 , buf_splittern279ton304n343_n304_6 );
buf_AQFP buf_splittern279ton304n343_n304_7_( clk_6 , buf_splittern279ton304n343_n304_6 , 0 , buf_splittern279ton304n343_n304_7 );
buf_AQFP buf_splittern279ton304n343_n304_8_( clk_8 , buf_splittern279ton304n343_n304_7 , 0 , buf_splittern279ton304n343_n304_8 );
buf_AQFP buf_splittern279ton304n343_n304_9_( clk_2 , buf_splittern279ton304n343_n304_8 , 0 , buf_splittern279ton304n343_n304_9 );
buf_AQFP buf_splittern279ton304n343_n337_1_( clk_2 , splittern279ton304n343 , 0 , buf_splittern279ton304n343_n337_1 );
buf_AQFP buf_splittern279ton304n343_n337_2_( clk_4 , buf_splittern279ton304n343_n337_1 , 0 , buf_splittern279ton304n343_n337_2 );
buf_AQFP buf_splittern279ton304n343_n337_3_( clk_6 , buf_splittern279ton304n343_n337_2 , 0 , buf_splittern279ton304n343_n337_3 );
buf_AQFP buf_splitterfromn280_n303_1_( clk_1 , splitterfromn280 , 0 , buf_splitterfromn280_n303_1 );
buf_AQFP buf_splitterfromn280_n303_2_( clk_3 , buf_splitterfromn280_n303_1 , 0 , buf_splitterfromn280_n303_2 );
buf_AQFP buf_splitterfromn280_n303_3_( clk_5 , buf_splitterfromn280_n303_2 , 0 , buf_splitterfromn280_n303_3 );
buf_AQFP buf_splitterfromn280_n303_4_( clk_7 , buf_splitterfromn280_n303_3 , 0 , buf_splitterfromn280_n303_4 );
buf_AQFP buf_splitterfromn280_n303_5_( clk_1 , buf_splitterfromn280_n303_4 , 0 , buf_splitterfromn280_n303_5 );
buf_AQFP buf_splittern287ton302n358_n302_1_( clk_2 , splittern287ton302n358 , 0 , buf_splittern287ton302n358_n302_1 );
buf_AQFP buf_splittern287ton302n358_n302_2_( clk_4 , buf_splittern287ton302n358_n302_1 , 0 , buf_splittern287ton302n358_n302_2 );
buf_AQFP buf_splittern287ton302n358_n302_3_( clk_6 , buf_splittern287ton302n358_n302_2 , 0 , buf_splittern287ton302n358_n302_3 );
buf_AQFP buf_splittern287ton302n358_n302_4_( clk_8 , buf_splittern287ton302n358_n302_3 , 0 , buf_splittern287ton302n358_n302_4 );
buf_AQFP buf_splittern287ton302n358_n302_5_( clk_2 , buf_splittern287ton302n358_n302_4 , 0 , buf_splittern287ton302n358_n302_5 );
buf_AQFP buf_splittern287ton302n358_n302_6_( clk_3 , buf_splittern287ton302n358_n302_5 , 0 , buf_splittern287ton302n358_n302_6 );
buf_AQFP buf_splittern287ton302n358_n302_7_( clk_4 , buf_splittern287ton302n358_n302_6 , 0 , buf_splittern287ton302n358_n302_7 );
buf_AQFP buf_splittern287ton302n358_n302_8_( clk_5 , buf_splittern287ton302n358_n302_7 , 0 , buf_splittern287ton302n358_n302_8 );
buf_AQFP buf_splittern287ton302n358_n302_9_( clk_7 , buf_splittern287ton302n358_n302_8 , 0 , buf_splittern287ton302n358_n302_9 );
buf_AQFP buf_splitterfromn288_n301_1_( clk_3 , splitterfromn288 , 0 , buf_splitterfromn288_n301_1 );
buf_AQFP buf_splitterfromn288_n301_2_( clk_5 , buf_splitterfromn288_n301_1 , 0 , buf_splitterfromn288_n301_2 );
buf_AQFP buf_splitterfromn288_n301_3_( clk_7 , buf_splitterfromn288_n301_2 , 0 , buf_splitterfromn288_n301_3 );
buf_AQFP buf_splitterfromn288_n301_4_( clk_1 , buf_splitterfromn288_n301_3 , 0 , buf_splitterfromn288_n301_4 );
buf_AQFP buf_splitterfromn288_n301_5_( clk_2 , buf_splitterfromn288_n301_4 , 0 , buf_splitterfromn288_n301_5 );
buf_AQFP buf_splitterfromn288_n301_6_( clk_3 , buf_splitterfromn288_n301_5 , 0 , buf_splitterfromn288_n301_6 );
buf_AQFP buf_splitterfromn288_n301_7_( clk_4 , buf_splitterfromn288_n301_6 , 0 , buf_splitterfromn288_n301_7 );
buf_AQFP buf_splitterfromn288_n301_8_( clk_6 , buf_splitterfromn288_n301_7 , 0 , buf_splitterfromn288_n301_8 );
buf_AQFP buf_splittern295ton300n313_n300_1_( clk_3 , splittern295ton300n313 , 0 , buf_splittern295ton300n313_n300_1 );
buf_AQFP buf_splittern295ton300n313_n300_2_( clk_5 , buf_splittern295ton300n313_n300_1 , 0 , buf_splittern295ton300n313_n300_2 );
buf_AQFP buf_splittern295ton300n313_n300_3_( clk_7 , buf_splittern295ton300n313_n300_2 , 0 , buf_splittern295ton300n313_n300_3 );
buf_AQFP buf_splittern295ton300n313_n300_4_( clk_1 , buf_splittern295ton300n313_n300_3 , 0 , buf_splittern295ton300n313_n300_4 );
buf_AQFP buf_splittern295ton300n313_n300_5_( clk_3 , buf_splittern295ton300n313_n300_4 , 0 , buf_splittern295ton300n313_n300_5 );
buf_AQFP buf_splittern295ton300n313_n300_6_( clk_4 , buf_splittern295ton300n313_n300_5 , 0 , buf_splittern295ton300n313_n300_6 );
buf_AQFP buf_splittern295ton300n313_n307_1_( clk_2 , splittern295ton300n313 , 0 , buf_splittern295ton300n313_n307_1 );
buf_AQFP buf_splitterfromn296_n299_1_( clk_3 , splitterfromn296 , 0 , buf_splitterfromn296_n299_1 );
buf_AQFP buf_splitterfromn296_n299_2_( clk_5 , buf_splitterfromn296_n299_1 , 0 , buf_splitterfromn296_n299_2 );
buf_AQFP buf_splitterfromn296_n299_3_( clk_7 , buf_splitterfromn296_n299_2 , 0 , buf_splitterfromn296_n299_3 );
buf_AQFP buf_splitterfromn296_n299_4_( clk_1 , buf_splitterfromn296_n299_3 , 0 , buf_splitterfromn296_n299_4 );
buf_AQFP buf_splitterfromn296_n299_5_( clk_3 , buf_splitterfromn296_n299_4 , 0 , buf_splitterfromn296_n299_5 );
buf_AQFP buf_splittern298ton299n312_n312_1_( clk_5 , splittern298ton299n312 , 0 , buf_splittern298ton299n312_n312_1 );
buf_AQFP buf_splitterfromn307_n310_1_( clk_2 , splitterfromn307 , 0 , buf_splitterfromn307_n310_1 );
buf_AQFP buf_splitterfromn307_n310_2_( clk_4 , buf_splitterfromn307_n310_1 , 0 , buf_splitterfromn307_n310_2 );
buf_AQFP buf_splitterfromn307_n310_3_( clk_6 , buf_splitterfromn307_n310_2 , 0 , buf_splitterfromn307_n310_3 );
buf_AQFP buf_splitterfromn307_n311_1_( clk_2 , splitterfromn307 , 0 , buf_splitterfromn307_n311_1 );
buf_AQFP buf_splitterfromn307_n311_2_( clk_4 , buf_splitterfromn307_n311_1 , 0 , buf_splitterfromn307_n311_2 );
buf_AQFP buf_splittern322ton323n327_n323_1_( clk_4 , splittern322ton323n327 , 0 , buf_splittern322ton323n327_n323_1 );
buf_AQFP buf_splittern322ton323n327_n323_2_( clk_6 , buf_splittern322ton323n327_n323_1 , 0 , buf_splittern322ton323n327_n323_2 );
buf_AQFP buf_splittern322ton323n327_n323_3_( clk_8 , buf_splittern322ton323n327_n323_2 , 0 , buf_splittern322ton323n327_n323_3 );
buf_AQFP buf_splittern322ton323n327_n323_4_( clk_2 , buf_splittern322ton323n327_n323_3 , 0 , buf_splittern322ton323n327_n323_4 );
buf_AQFP buf_splittern322ton323n327_n323_5_( clk_4 , buf_splittern322ton323n327_n323_4 , 0 , buf_splittern322ton323n327_n323_5 );
buf_AQFP buf_splittern322ton323n327_n323_6_( clk_6 , buf_splittern322ton323n327_n323_5 , 0 , buf_splittern322ton323n327_n323_6 );
buf_AQFP buf_splittern322ton323n327_n323_7_( clk_8 , buf_splittern322ton323n327_n323_6 , 0 , buf_splittern322ton323n327_n323_7 );
buf_AQFP buf_splittern322ton323n327_n323_8_( clk_2 , buf_splittern322ton323n327_n323_7 , 0 , buf_splittern322ton323n327_n323_8 );
buf_AQFP buf_splittern322ton323n327_n323_9_( clk_4 , buf_splittern322ton323n327_n323_8 , 0 , buf_splittern322ton323n327_n323_9 );
buf_AQFP buf_splittern322ton323n327_n324_1_( clk_4 , splittern322ton323n327 , 0 , buf_splittern322ton323n327_n324_1 );
buf_AQFP buf_splittern322ton323n327_n324_2_( clk_6 , buf_splittern322ton323n327_n324_1 , 0 , buf_splittern322ton323n327_n324_2 );
buf_AQFP buf_splittern322ton323n327_n324_3_( clk_8 , buf_splittern322ton323n327_n324_2 , 0 , buf_splittern322ton323n327_n324_3 );
buf_AQFP buf_splittern322ton323n327_n324_4_( clk_2 , buf_splittern322ton323n327_n324_3 , 0 , buf_splittern322ton323n327_n324_4 );
buf_AQFP buf_splittern322ton323n327_n324_5_( clk_4 , buf_splittern322ton323n327_n324_4 , 0 , buf_splittern322ton323n327_n324_5 );
buf_AQFP buf_splittern322ton323n327_n324_6_( clk_6 , buf_splittern322ton323n327_n324_5 , 0 , buf_splittern322ton323n327_n324_6 );
buf_AQFP buf_splittern322ton323n327_n324_7_( clk_8 , buf_splittern322ton323n327_n324_6 , 0 , buf_splittern322ton323n327_n324_7 );
buf_AQFP buf_splittern322ton323n327_n324_8_( clk_2 , buf_splittern322ton323n327_n324_7 , 0 , buf_splittern322ton323n327_n324_8 );
buf_AQFP buf_splittern322ton323n327_n324_9_( clk_4 , buf_splittern322ton323n327_n324_8 , 0 , buf_splittern322ton323n327_n324_9 );
buf_AQFP buf_splittern322ton323n327_n324_10_( clk_6 , buf_splittern322ton323n327_n324_9 , 0 , buf_splittern322ton323n327_n324_10 );
buf_AQFP buf_splittern337ton338n342_n338_1_( clk_8 , splittern337ton338n342 , 0 , buf_splittern337ton338n342_n338_1 );
buf_AQFP buf_splittern337ton338n342_n338_2_( clk_2 , buf_splittern337ton338n342_n338_1 , 0 , buf_splittern337ton338n342_n338_2 );
buf_AQFP buf_splittern337ton338n342_n338_3_( clk_3 , buf_splittern337ton338n342_n338_2 , 0 , buf_splittern337ton338n342_n338_3 );
buf_AQFP buf_splittern337ton338n342_n339_1_( clk_7 , splittern337ton338n342 , 0 , buf_splittern337ton338n342_n339_1 );
buf_AQFP buf_splittern337ton338n342_n339_2_( clk_8 , buf_splittern337ton338n342_n339_1 , 0 , buf_splittern337ton338n342_n339_2 );
buf_AQFP buf_splittern337ton338n342_n339_3_( clk_1 , buf_splittern337ton338n342_n339_2 , 0 , buf_splittern337ton338n342_n339_3 );
buf_AQFP buf_splittern337ton338n342_n339_4_( clk_2 , buf_splittern337ton338n342_n339_3 , 0 , buf_splittern337ton338n342_n339_4 );
buf_AQFP buf_splittern337ton338n342_n339_5_( clk_3 , buf_splittern337ton338n342_n339_4 , 0 , buf_splittern337ton338n342_n339_5 );
buf_AQFP buf_splittern352ton353n357_n353_1_( clk_5 , splittern352ton353n357 , 0 , buf_splittern352ton353n357_n353_1 );
buf_AQFP buf_splittern352ton353n357_n353_2_( clk_6 , buf_splittern352ton353n357_n353_1 , 0 , buf_splittern352ton353n357_n353_2 );
buf_AQFP buf_splittern352ton353n357_n353_3_( clk_7 , buf_splittern352ton353n357_n353_2 , 0 , buf_splittern352ton353n357_n353_3 );
buf_AQFP buf_splittern352ton353n357_n353_4_( clk_8 , buf_splittern352ton353n357_n353_3 , 0 , buf_splittern352ton353n357_n353_4 );
buf_AQFP buf_splittern352ton353n357_n353_5_( clk_2 , buf_splittern352ton353n357_n353_4 , 0 , buf_splittern352ton353n357_n353_5 );
buf_AQFP buf_splittern352ton353n357_n353_6_( clk_4 , buf_splittern352ton353n357_n353_5 , 0 , buf_splittern352ton353n357_n353_6 );
buf_AQFP buf_splittern352ton353n357_n353_7_( clk_6 , buf_splittern352ton353n357_n353_6 , 0 , buf_splittern352ton353n357_n353_7 );
buf_AQFP buf_splittern352ton353n357_n354_1_( clk_6 , splittern352ton353n357 , 0 , buf_splittern352ton353n357_n354_1 );
buf_AQFP buf_splittern352ton353n357_n354_2_( clk_8 , buf_splittern352ton353n357_n354_1 , 0 , buf_splittern352ton353n357_n354_2 );
buf_AQFP buf_splittern352ton353n357_n354_3_( clk_2 , buf_splittern352ton353n357_n354_2 , 0 , buf_splittern352ton353n357_n354_3 );
buf_AQFP buf_splittern352ton353n357_n354_4_( clk_4 , buf_splittern352ton353n357_n354_3 , 0 , buf_splittern352ton353n357_n354_4 );
buf_AQFP buf_splittern352ton353n357_n354_5_( clk_6 , buf_splittern352ton353n357_n354_4 , 0 , buf_splittern352ton353n357_n354_5 );
buf_AQFP buf_splittern352ton353n357_n354_6_( clk_7 , buf_splittern352ton353n357_n354_5 , 0 , buf_splittern352ton353n357_n354_6 );
splitter_AQFP splitterN1ton147n70_( clk_2 , N1 , 0 , splitterN1ton147n70 );
splitter_AQFP splitterN101ton102n316_( clk_4 , buf_N101_splitterN101ton102n316_1 , 0 , splitterN101ton102n316 );
splitter_AQFP splitterN106ton102n289_( clk_5 , buf_N106_splitterN106ton102n289_1 , 0 , splitterN106ton102n289 );
splitter_AQFP splitterN111ton105n237_( clk_5 , buf_N111_splitterN111ton105n237_1 , 0 , splitterN111ton105n237 );
splitter_AQFP splitterN116ton105n255_( clk_5 , buf_N116_splitterN116ton105n255_1 , 0 , splitterN116ton105n255 );
splitter_AQFP splitterN121ton182n97_( clk_5 , buf_N121_splitterN121ton182n97_2 , 0 , splitterN121ton182n97 );
splitter_AQFP splitterN126ton100n99_( clk_7 , buf_N126_splitterN126ton100n99_2 , 0 , splitterN126ton100n99 );
splitter_AQFP splitterfromN13_( clk_5 , buf_N13_splitterfromN13_1 , 0 , splitterfromN13 );
splitter_AQFP splitterN130ton120n91_( clk_2 , N130 , 0 , splitterN130ton120n91 );
splitter_AQFP splitterfromN135_( clk_4 , buf_N135_splitterfromN135_1 , 0 , splitterfromN135 );
splitter_AQFP splitterN138ton267n291_( clk_7 , buf_N138_splitterN138ton267n291_2 , 0 , splitterN138ton267n291 );
splitter_AQFP splitterfromN143_( clk_2 , buf_N143_splitterfromN143_5 , 0 , splitterfromN143 );
splitter_AQFP splitterfromN146_( clk_7 , buf_N146_splitterfromN146_2 , 0 , splitterfromN146 );
splitter_AQFP splitterfromN149_( clk_2 , buf_N149_splitterfromN149_4 , 0 , splitterfromN149 );
splitter_AQFP splitterfromN153_( clk_6 , buf_N153_splitterfromN153_2 , 0 , splitterfromN153 );
splitter_AQFP splitterN159ton117n330_( clk_4 , buf_N159_splitterN159ton117n330_1 , 0 , splitterN159ton117n330 );
splitter_AQFP splitterN159ton272n330_( clk_5 , splitterN159ton117n330 , 0 , splitterN159ton272n330 );
splitter_AQFP splitterN165ton129n346_( clk_6 , buf_N165_splitterN165ton129n346_2 , 0 , splitterN165ton129n346 );
splitter_AQFP splitterN165ton280n346_( clk_5 , splitterN165ton129n346 , 0 , splitterN165ton280n346 );
splitter_AQFP splitterN17ton146n68_( clk_2 , N17 , 0 , splitterN17ton146n68 );
splitter_AQFP splitterN17ton159n68_( clk_3 , splitterN17ton146n68 , 0 , splitterN17ton159n68 );
splitter_AQFP splitterN171ton132n361_( clk_8 , buf_N171_splitterN171ton132n361_3 , 0 , splitterN171ton132n361 );
splitter_AQFP splitterN171ton288n361_( clk_4 , splitterN171ton132n361 , 0 , splitterN171ton288n361 );
splitter_AQFP splitterN177ton117n315_( clk_5 , buf_N177_splitterN177ton117n315_2 , 0 , splitterN177ton117n315 );
splitter_AQFP splitterN177ton296n315_( clk_4 , splitterN177ton117n315 , 0 , splitterN177ton296n315 );
splitter_AQFP splitterN183ton132n221_( clk_8 , buf_N183_splitterN183ton132n221_3 , 0 , splitterN183ton132n221 );
splitter_AQFP splitterN183ton212n221_( clk_3 , splitterN183ton132n221 , 0 , splitterN183ton212n221 );
splitter_AQFP splitterN189ton123n236_( clk_5 , buf_N189_splitterN189ton123n236_1 , 0 , splitterN189ton123n236 );
splitter_AQFP splitterN189ton194n236_( clk_5 , splitterN189ton123n236 , 0 , splitterN189ton194n236 );
splitter_AQFP splitterN195ton123n253_( clk_8 , buf_N195_splitterN195ton123n253_4 , 0 , splitterN195ton123n253 );
splitter_AQFP splitterN195ton200n253_( clk_4 , splitterN195ton123n253 , 0 , splitterN195ton200n253 );
splitter_AQFP splitterN201ton129n180_( clk_5 , buf_N201_splitterN201ton129n180_1 , 0 , splitterN201ton129n180 );
splitter_AQFP splitterN201ton167n180_( clk_3 , splitterN201ton129n180 , 0 , splitterN201ton167n180 );
splitter_AQFP splitterfromN207_( clk_3 , buf_N207_splitterfromN207_6 , 0 , splitterfromN207 );
splitter_AQFP splitterN210ton182n360_( clk_5 , buf_N210_splitterN210ton182n360_1 , 0 , splitterN210ton182n360 );
splitter_AQFP splitterN210ton237n255_( clk_6 , splitterN210ton182n360 , 0 , splitterN210ton237n255 );
splitter_AQFP splitterN210ton316n360_( clk_7 , splitterN210ton182n360 , 0 , splitterN210ton316n360 );
splitter_AQFP splitterN219ton171n355_( clk_5 , buf_N219_splitterN219ton171n355_5 , 0 , splitterN219ton171n355 );
splitter_AQFP splitterN219ton232n308_( clk_5 , splitterN219ton171n355 , 0 , splitterN219ton232n308 );
splitter_AQFP splitterN219ton311n355_( clk_5 , splitterN219ton171n355 , 0 , splitterN219ton311n355 );
splitter_AQFP splitterN228ton173n357_( clk_7 , buf_N228_splitterN228ton173n357_8 , 0 , splitterN228ton173n357 );
splitter_AQFP splitterN228ton233n250_( clk_2 , splitterN228ton173n357 , 0 , splitterN228ton233n250 );
splitter_AQFP splitterN228ton309n357_( clk_4 , splitterN228ton173n357 , 0 , splitterN228ton309n357 );
splitter_AQFP splitterN237ton174n358_( clk_5 , buf_N237_splitterN237ton174n358_1 , 0 , splitterN237ton174n358 );
splitter_AQFP splitterN237ton234n251_( clk_8 , splitterN237ton174n358 , 0 , splitterN237ton234n251 );
splitter_AQFP splitterN237ton313n358_( clk_6 , splitterN237ton174n358 , 0 , splitterN237ton313n358 );
splitter_AQFP splitterN246ton175n359_( clk_4 , buf_N246_splitterN246ton175n359_5 , 0 , splitterN246ton175n359 );
splitter_AQFP splitterN246ton235n252_( clk_6 , splitterN246ton175n359 , 0 , splitterN246ton235n252 );
splitter_AQFP splitterN246ton314n359_( clk_5 , splitterN246ton175n359 , 0 , splitterN246ton314n359 );
splitter_AQFP splitterN255ton181n254_( clk_5 , buf_N255_splitterN255ton181n254_1 , 0 , splitterN255ton181n254 );
splitter_AQFP splitterN261ton169n201_( clk_3 , buf_N261_splitterN261ton169n201_4 , 0 , splitterN261ton169n201 );
splitter_AQFP splitterN268ton152n331_( clk_4 , buf_N268_splitterN268ton152n331_1 , 0 , splitterN268ton152n331 );
splitter_AQFP splitterN29ton61n84_( clk_2 , N29 , 0 , splitterN29ton61n84 );
splitter_AQFP splitterfromN36_( clk_2 , N36 , 0 , splitterfromN36 );
splitter_AQFP splitterN42ton153n77_( clk_3 , N42 , 0 , splitterN42ton153n77 );
splitter_AQFP splitterN42ton176n77_( clk_5 , splitterN42ton153n77 , 0 , splitterN42ton176n77 );
splitter_AQFP splitterN51ton159n81_( clk_4 , buf_N51_splitterN51ton159n81_1 , 0 , splitterN51ton159n81 );
splitter_AQFP splitterN55ton151n82_( clk_5 , buf_N55_splitterN55ton151n82_2 , 0 , splitterN55ton151n82 );
splitter_AQFP splitterN59ton144n86_( clk_2 , N59 , 0 , splitterN59ton144n86 );
splitter_AQFP splitterfromN68_( clk_3 , N68 , 0 , splitterfromN68 );
splitter_AQFP splitterfromN75_( clk_2 , N75 , 0 , splitterfromN75 );
splitter_AQFP splitterfromN8_( clk_2 , N8 , 0 , splitterfromN8 );
splitter_AQFP splitterN80ton149n76_( clk_5 , buf_N80_splitterN80ton149n76_2 , 0 , splitterN80ton149n76 );
splitter_AQFP splitterN91ton262n94_( clk_6 , buf_N91_splitterN91ton262n94_2 , 0 , splitterN91ton262n94 );
splitter_AQFP splitterN96ton273n91_( clk_3 , N96 , 0 , splitterN96ton273n91 );
splitter_AQFP splitterfromn61_( clk_5 , n61 , 0 , splitterfromn61 );
splitter_AQFP splitterfromn63_( clk_8 , buf_n63_splitterfromn63_2 , 0 , splitterfromn63 );
splitter_AQFP splittern65toN390n80_( clk_2 , buf_n65_splittern65toN390n80_15 , 0 , splittern65toN390n80 );
splitter_AQFP splittern67ton160n83_( clk_6 , buf_n67_splittern67ton160n83_1 , 0 , splittern67ton160n83 );
splitter_AQFP splitterfromn68_( clk_1 , buf_n68_splitterfromn68_4 , 0 , splitterfromn68 );
splitter_AQFP splitterfromn70_( clk_4 , n70 , 0 , splitterfromn70 );
splitter_AQFP splitterfromn71_( clk_7 , buf_n71_splitterfromn71_5 , 0 , splitterfromn71 );
splitter_AQFP splitterfromn73_( clk_6 , buf_n73_splitterfromn73_1 , 0 , splitterfromn73 );
splitter_AQFP splitterfromn75_( clk_4 , n75 , 0 , splitterfromn75 );
splitter_AQFP splitterfromn78_( clk_4 , n78 , 0 , splitterfromn78 );
splitter_AQFP splittern81toN447n156_( clk_6 , n81 , 0 , splittern81toN447n156 );
splitter_AQFP splittern83ton179n88_( clk_1 , n83 , 0 , splittern83ton179n88 );
splitter_AQFP splitterfromn86_( clk_6 , n86 , 0 , splitterfromn86 );
splitter_AQFP splitterfromn92_( clk_6 , n92 , 0 , splitterfromn92 );
splitter_AQFP splitterfromn95_( clk_3 , buf_n95_splitterfromn95_3 , 0 , splitterfromn95 );
splitter_AQFP splitterfromn98_( clk_8 , n98 , 0 , splitterfromn98 );
splitter_AQFP splitterfromn101_( clk_4 , n101 , 0 , splitterfromn101 );
splitter_AQFP splitterfromn104_( clk_8 , n104 , 0 , splitterfromn104 );
splitter_AQFP splitterfromn107_( clk_1 , n107 , 0 , splitterfromn107 );
splitter_AQFP splitterfromn110_( clk_5 , n110 , 0 , splitterfromn110 );
splitter_AQFP splitterfromn113_( clk_6 , buf_n113_splitterfromn113_2 , 0 , splitterfromn113 );
splitter_AQFP splitterfromn119_( clk_3 , buf_n119_splitterfromn119_1 , 0 , splitterfromn119 );
splitter_AQFP splitterfromn122_( clk_6 , buf_n122_splitterfromn122_3 , 0 , splitterfromn122 );
splitter_AQFP splitterfromn125_( clk_4 , n125 , 0 , splitterfromn125 );
splitter_AQFP splitterfromn128_( clk_8 , n128 , 0 , splitterfromn128 );
splitter_AQFP splitterfromn131_( clk_3 , n131 , 0 , splitterfromn131 );
splitter_AQFP splitterfromn134_( clk_3 , n134 , 0 , splitterfromn134 );
splitter_AQFP splitterfromn137_( clk_1 , n137 , 0 , splitterfromn137 );
splitter_AQFP splitterfromn140_( clk_1 , buf_n140_splitterfromn140_2 , 0 , splitterfromn140 );
splitter_AQFP splitterfromn144_( clk_4 , n144 , 0 , splitterfromn144 );
splitter_AQFP splitterfromn145_( clk_8 , n145 , 0 , splitterfromn145 );
splitter_AQFP splittern147ton148n208_( clk_3 , n147 , 0 , splittern147ton148n208 );
splitter_AQFP splitterfromn150_( clk_8 , n150 , 0 , splitterfromn150 );
splitter_AQFP splittern152ton164n210_( clk_3 , n152 , 0 , splittern152ton164n210 );
splitter_AQFP splittern162ton163n289_( clk_2 , n162 , 0 , splittern162ton163n289 );
splitter_AQFP splittern162ton196n207_( clk_3 , splittern162ton163n289 , 0 , splittern162ton196n207 );
splitter_AQFP splittern162ton262n289_( clk_3 , splittern162ton163n289 , 0 , splittern162ton262n289 );
splitter_AQFP splittern165ton166n175_( clk_6 , n165 , 0 , splittern165ton166n175 );
splitter_AQFP splitterfromn166_( clk_8 , n166 , 0 , splitterfromn166 );
splitter_AQFP splittern167ton168n201_( clk_8 , n167 , 0 , splittern167ton168n201 );
splitter_AQFP splittern168ton169n173_( clk_2 , n168 , 0 , splittern168ton169n173 );
splitter_AQFP splittern179ton180n361_( clk_3 , n179 , 0 , splittern179ton180n361 );
splitter_AQFP splittern179ton236n253_( clk_5 , splittern179ton180n361 , 0 , splittern179ton236n253 );
splitter_AQFP splittern179ton315n361_( clk_4 , splittern179ton180n361 , 0 , splittern179ton315n361 );
splitter_AQFP splittern192ton193n235_( clk_6 , n192 , 0 , splittern192ton193n235 );
splitter_AQFP splittern193ton206n234_( clk_8 , n193 , 0 , splittern193ton206n234 );
splitter_AQFP splitterfromn194_( clk_8 , n194 , 0 , splitterfromn194 );
splitter_AQFP splittern198ton199n252_( clk_7 , n198 , 0 , splittern198ton199n252 );
splitter_AQFP splittern199ton204n251_( clk_1 , n199 , 0 , splittern199ton204n251 );
splitter_AQFP splitterfromn200_( clk_1 , n200 , 0 , splitterfromn200 );
splitter_AQFP splittern202ton203n247_( clk_3 , n202 , 0 , splittern202ton203n247 );
splitter_AQFP splittern204ton205n230_( clk_6 , n204 , 0 , splittern204ton205n230 );
splitter_AQFP splittern206ton214n297_( clk_1 , n206 , 0 , splittern206ton214n297 );
splitter_AQFP splittern210ton211n220_( clk_7 , n210 , 0 , splittern210ton211n220 );
splitter_AQFP splittern211ton213n298_( clk_1 , n211 , 0 , splittern211ton213n298 );
splitter_AQFP splitterfromn212_( clk_1 , n212 , 0 , splitterfromn212 );
splitter_AQFP splittern213ton214n218_( clk_3 , n213 , 0 , splittern213ton214n218 );
splitter_AQFP splittern228ton229n233_( clk_2 , n228 , 0 , splittern228ton229n233 );
splitter_AQFP splittern245ton246n250_( clk_3 , n245 , 0 , splittern245ton246n250 );
splitter_AQFP splittern263ton264n290_( clk_2 , n263 , 0 , splittern263ton264n290 );
splitter_AQFP splittern266ton268n292_( clk_2 , n266 , 0 , splittern266ton268n292 );
splitter_AQFP splittern270ton271n329_( clk_6 , n270 , 0 , splittern270ton271n329 );
splitter_AQFP splittern271ton306n328_( clk_8 , n271 , 0 , splittern271ton306n328 );
splitter_AQFP splitterfromn272_( clk_1 , n272 , 0 , splitterfromn272 );
splitter_AQFP splittern278ton279n344_( clk_6 , n278 , 0 , splittern278ton279n344 );
splitter_AQFP splittern279ton304n343_( clk_8 , n279 , 0 , splittern279ton304n343 );
splitter_AQFP splitterfromn280_( clk_7 , buf_n280_splitterfromn280_4 , 0 , splitterfromn280 );
splitter_AQFP splittern286ton287n359_( clk_6 , n286 , 0 , splittern286ton287n359 );
splitter_AQFP splittern287ton302n358_( clk_8 , n287 , 0 , splittern287ton302n358 );
splitter_AQFP splitterfromn288_( clk_1 , n288 , 0 , splitterfromn288 );
splitter_AQFP splittern294ton295n314_( clk_6 , n294 , 0 , splittern294ton295n314 );
splitter_AQFP splittern295ton300n313_( clk_1 , n295 , 0 , splittern295ton300n313 );
splitter_AQFP splitterfromn296_( clk_2 , n296 , 0 , splitterfromn296 );
splitter_AQFP splittern298ton299n312_( clk_4 , n298 , 0 , splittern298ton299n312 );
splitter_AQFP splittern300ton301n354_( clk_7 , n300 , 0 , splittern300ton301n354 );
splitter_AQFP splittern302ton303n339_( clk_2 , n302 , 0 , splittern302ton303n339 );
splitter_AQFP splittern304ton305n324_( clk_5 , n304 , 0 , splittern304ton305n324 );
splitter_AQFP splitterfromn307_( clk_8 , buf_n307_splitterfromn307_1 , 0 , splitterfromn307 );
splitter_AQFP splittern322ton323n327_( clk_3 , n322 , 0 , splittern322ton323n327 );
splitter_AQFP splittern337ton338n342_( clk_6 , buf_n337_splittern337ton338n342_3 , 0 , splittern337ton338n342 );
splitter_AQFP splittern352ton353n357_( clk_4 , n352 , 0 , splittern352ton353n357 );

endmodule