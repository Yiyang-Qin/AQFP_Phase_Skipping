module top( clk_1 , clk_2 , clk_3 , clk_4 , clk_5 , clk_6 , clk_7 , clk_8 , N1 , N102 , N105 , N108 , N11 , N112 , N115 , N14 , N17 , N21 , N24 , N27 , N30 , N34 , N37 , N4 , N40 , N43 , N47 , N50 , N53 , N56 , N60 , N63 , N66 , N69 , N73 , N76 , N79 , N8 , N82 , N86 , N89 , N92 , N95 , N99 , N223 , N329 , N370 , N421 , N430 , N431 , N432 );

input N1 , N102 , N105 , N108 , N11 , N112 , N115 , N14 , N17 , N21 , N24 , N27 , N30 , N34 , N37 , N4 , N40 , N43 , N47 , N50 , N53 , N56 , N60 , N63 , N66 , N69 , N73 , N76 , N79 , N8 , N82 , N86 , N89 , N92 , N95 , N99 ;
output N223 , N329 , N370 , N421 , N430 , N431 , N432 ;
wire n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , buf_N102_splitterfromN102_1 , buf_N105_splitterfromN105_10 , buf_N105_splitterfromN105_9 , buf_N105_splitterfromN105_8 , buf_N105_splitterfromN105_7 , buf_N105_splitterfromN105_6 , buf_N105_splitterfromN105_5 , buf_N105_splitterfromN105_4 , buf_N105_splitterfromN105_3 , buf_N105_splitterfromN105_2 , buf_N105_splitterfromN105_1 , buf_N108_splitterfromN108_1 , buf_N112_splitterfromN112_5 , buf_N112_splitterfromN112_4 , buf_N112_splitterfromN112_3 , buf_N112_splitterfromN112_2 , buf_N112_splitterfromN112_1 , buf_N115_splitterfromN115_10 , buf_N115_splitterfromN115_9 , buf_N115_splitterfromN115_8 , buf_N115_splitterfromN115_7 , buf_N115_splitterfromN115_6 , buf_N115_splitterfromN115_5 , buf_N115_splitterfromN115_4 , buf_N115_splitterfromN115_3 , buf_N115_splitterfromN115_2 , buf_N115_splitterfromN115_1 , buf_N14_splitterfromN14_10 , buf_N14_splitterfromN14_9 , buf_N14_splitterfromN14_8 , buf_N14_splitterfromN14_7 , buf_N14_splitterfromN14_6 , buf_N14_splitterfromN14_5 , buf_N14_splitterfromN14_4 , buf_N14_splitterfromN14_3 , buf_N14_splitterfromN14_2 , buf_N14_splitterfromN14_1 , buf_N21_splitterfromN21_5 , buf_N21_splitterfromN21_4 , buf_N21_splitterfromN21_3 , buf_N21_splitterfromN21_2 , buf_N21_splitterfromN21_1 , buf_N24_n37_1 , buf_N27_splitterfromN27_10 , buf_N27_splitterfromN27_9 , buf_N27_splitterfromN27_8 , buf_N27_splitterfromN27_7 , buf_N27_splitterfromN27_6 , buf_N27_splitterfromN27_5 , buf_N27_splitterfromN27_4 , buf_N27_splitterfromN27_3 , buf_N27_splitterfromN27_2 , buf_N27_splitterfromN27_1 , buf_N34_splitterfromN34_5 , buf_N34_splitterfromN34_4 , buf_N34_splitterfromN34_3 , buf_N34_splitterfromN34_2 , buf_N34_splitterfromN34_1 , buf_N4_splitterfromN4_1 , buf_N40_splitterfromN40_10 , buf_N40_splitterfromN40_9 , buf_N40_splitterfromN40_8 , buf_N40_splitterfromN40_7 , buf_N40_splitterfromN40_6 , buf_N40_splitterfromN40_5 , buf_N40_splitterfromN40_4 , buf_N40_splitterfromN40_3 , buf_N40_splitterfromN40_2 , buf_N40_splitterfromN40_1 , buf_N47_splitterfromN47_5 , buf_N47_splitterfromN47_4 , buf_N47_splitterfromN47_3 , buf_N47_splitterfromN47_2 , buf_N47_splitterfromN47_1 , buf_N53_splitterfromN53_10 , buf_N53_splitterfromN53_9 , buf_N53_splitterfromN53_8 , buf_N53_splitterfromN53_7 , buf_N53_splitterfromN53_6 , buf_N53_splitterfromN53_5 , buf_N53_splitterfromN53_4 , buf_N53_splitterfromN53_3 , buf_N53_splitterfromN53_2 , buf_N53_splitterfromN53_1 , buf_N60_splitterfromN60_5 , buf_N60_splitterfromN60_4 , buf_N60_splitterfromN60_3 , buf_N60_splitterfromN60_2 , buf_N60_splitterfromN60_1 , buf_N66_n112_10 , buf_N66_n112_9 , buf_N66_n112_8 , buf_N66_n112_7 , buf_N66_n112_6 , buf_N66_n112_5 , buf_N66_n112_4 , buf_N66_n112_3 , buf_N66_n112_2 , buf_N66_n112_1 , buf_N73_splitterfromN73_5 , buf_N73_splitterfromN73_4 , buf_N73_splitterfromN73_3 , buf_N73_splitterfromN73_2 , buf_N73_splitterfromN73_1 , buf_N79_splitterfromN79_10 , buf_N79_splitterfromN79_9 , buf_N79_splitterfromN79_8 , buf_N79_splitterfromN79_7 , buf_N79_splitterfromN79_6 , buf_N79_splitterfromN79_5 , buf_N79_splitterfromN79_4 , buf_N79_splitterfromN79_3 , buf_N79_splitterfromN79_2 , buf_N79_splitterfromN79_1 , buf_N8_splitterfromN8_5 , buf_N8_splitterfromN8_4 , buf_N8_splitterfromN8_3 , buf_N8_splitterfromN8_2 , buf_N8_splitterfromN8_1 , buf_N86_splitterfromN86_5 , buf_N86_splitterfromN86_4 , buf_N86_splitterfromN86_3 , buf_N86_splitterfromN86_2 , buf_N86_splitterfromN86_1 , buf_N92_splitterfromN92_10 , buf_N92_splitterfromN92_9 , buf_N92_splitterfromN92_8 , buf_N92_splitterfromN92_7 , buf_N92_splitterfromN92_6 , buf_N92_splitterfromN92_5 , buf_N92_splitterfromN92_4 , buf_N92_splitterfromN92_3 , buf_N92_splitterfromN92_2 , buf_N92_splitterfromN92_1 , buf_N99_splitterfromN99_5 , buf_N99_splitterfromN99_4 , buf_N99_splitterfromN99_3 , buf_N99_splitterfromN99_2 , buf_N99_splitterfromN99_1 , buf_n148_n149_2 , buf_n148_n149_1 , buf_n151_N431_1 , buf_splitterfromN1_n69_3 , buf_splitterfromN1_n69_2 , buf_splitterfromN1_n69_1 , buf_splitterfromN102_n54_2 , buf_splitterfromN102_n54_1 , buf_splitterfromN105_n140_3 , buf_splitterfromN105_n140_2 , buf_splitterfromN105_n140_1 , buf_splitterfromN108_n55_3 , buf_splitterfromN108_n55_2 , buf_splitterfromN108_n55_1 , buf_splitterfromN11_n64_3 , buf_splitterfromN11_n64_2 , buf_splitterfromN11_n64_1 , buf_splitterfromN112_n117_3 , buf_splitterfromN112_n117_2 , buf_splitterfromN112_n117_1 , buf_splitterfromN115_n142_3 , buf_splitterfromN115_n142_2 , buf_splitterfromN115_n142_1 , buf_splitterfromN14_n147_3 , buf_splitterfromN14_n147_2 , buf_splitterfromN14_n147_1 , buf_splitterfromN17_n65_4 , buf_splitterfromN17_n65_3 , buf_splitterfromN17_n65_2 , buf_splitterfromN17_n65_1 , buf_splitterfromN21_n95_3 , buf_splitterfromN21_n95_2 , buf_splitterfromN21_n95_1 , buf_splitterfromN27_n126_2 , buf_splitterfromN27_n126_1 , buf_splitterfromN30_n61_3 , buf_splitterfromN30_n61_2 , buf_splitterfromN30_n61_1 , buf_splitterfromN34_n89_3 , buf_splitterfromN34_n89_2 , buf_splitterfromN34_n89_1 , buf_splitterfromN37_n82_3 , buf_splitterfromN37_n82_2 , buf_splitterfromN37_n82_1 , buf_splitterfromN4_n70_3 , buf_splitterfromN4_n70_2 , buf_splitterfromN4_n70_1 , buf_splitterfromN40_n124_2 , buf_splitterfromN40_n124_1 , buf_splitterfromN43_n83_3 , buf_splitterfromN43_n83_2 , buf_splitterfromN43_n83_1 , buf_splitterfromN47_n114_3 , buf_splitterfromN47_n114_2 , buf_splitterfromN47_n114_1 , buf_splitterfromN50_n76_3 , buf_splitterfromN50_n76_2 , buf_splitterfromN50_n76_1 , buf_splitterfromN53_n129_3 , buf_splitterfromN53_n129_2 , buf_splitterfromN53_n129_1 , buf_splitterfromN56_n77_4 , buf_splitterfromN56_n77_3 , buf_splitterfromN56_n77_2 , buf_splitterfromN56_n77_1 , buf_splitterfromN60_n110_3 , buf_splitterfromN60_n110_2 , buf_splitterfromN60_n110_1 , buf_splitterfromN69_n79_3 , buf_splitterfromN69_n79_2 , buf_splitterfromN69_n79_1 , buf_splitterfromN73_n107_3 , buf_splitterfromN73_n107_2 , buf_splitterfromN73_n107_1 , buf_splitterfromN76_n57_3 , buf_splitterfromN76_n57_2 , buf_splitterfromN76_n57_1 , buf_splitterfromN79_n137_3 , buf_splitterfromN79_n137_2 , buf_splitterfromN79_n137_1 , buf_splitterfromN8_n100_3 , buf_splitterfromN8_n100_2 , buf_splitterfromN8_n100_1 , buf_splitterfromN82_n58_4 , buf_splitterfromN82_n58_3 , buf_splitterfromN82_n58_2 , buf_splitterfromN82_n58_1 , buf_splitterfromN86_n103_3 , buf_splitterfromN86_n103_2 , buf_splitterfromN86_n103_1 , buf_splitterfromN89_n72_3 , buf_splitterfromN89_n72_2 , buf_splitterfromN89_n72_1 , buf_splitterfromN92_n135_3 , buf_splitterfromN92_n135_2 , buf_splitterfromN92_n135_1 , buf_splitterfromN95_n73_4 , buf_splitterfromN95_n73_3 , buf_splitterfromN95_n73_2 , buf_splitterfromN95_n73_1 , buf_splitterfromN99_n92_2 , buf_splitterfromN99_n92_1 , buf_splitterfromn37_n62_2 , buf_splitterfromn37_n62_1 , buf_splitterfromn45_n80_3 , buf_splitterfromn45_n80_2 , buf_splitterfromn45_n80_1 , buf_splittern53ton69N223_N223_14 , buf_splittern53ton69N223_N223_13 , buf_splittern53ton69N223_N223_12 , buf_splittern53ton69N223_N223_11 , buf_splittern53ton69N223_N223_10 , buf_splittern53ton69N223_N223_9 , buf_splittern53ton69N223_N223_8 , buf_splittern53ton69N223_N223_7 , buf_splittern53ton69N223_N223_6 , buf_splittern53ton69N223_N223_5 , buf_splittern53ton69N223_N223_4 , buf_splittern53ton69N223_N223_3 , buf_splittern53ton69N223_N223_2 , buf_splittern53ton69N223_N223_1 , buf_splitterfromn55_n118_3 , buf_splitterfromn55_n118_2 , buf_splitterfromn55_n118_1 , buf_splitterfromn58_n104_3 , buf_splitterfromn58_n104_2 , buf_splitterfromn58_n104_1 , buf_splitterfromn62_n90_3 , buf_splitterfromn62_n90_2 , buf_splitterfromn62_n90_1 , buf_splitterfromn65_n96_3 , buf_splitterfromn65_n96_2 , buf_splitterfromn65_n96_1 , buf_splitterfromn70_n101_3 , buf_splitterfromn70_n101_2 , buf_splitterfromn70_n101_1 , buf_splitterfromn73_n93_3 , buf_splitterfromn73_n93_2 , buf_splitterfromn73_n93_1 , buf_splitterfromn77_n111_3 , buf_splitterfromn77_n111_2 , buf_splitterfromn77_n111_1 , buf_splitterfromn80_n108_4 , buf_splitterfromn80_n108_3 , buf_splitterfromn80_n108_2 , buf_splitterfromn80_n108_1 , buf_splitterfromn83_n115_4 , buf_splitterfromn83_n115_3 , buf_splitterfromn83_n115_2 , buf_splitterfromn83_n115_1 , buf_splittern88ton117N329_N329_9 , buf_splittern88ton117N329_N329_8 , buf_splittern88ton117N329_N329_7 , buf_splittern88ton117N329_N329_6 , buf_splittern88ton117N329_N329_5 , buf_splittern88ton117N329_N329_4 , buf_splittern88ton117N329_N329_3 , buf_splittern88ton117N329_N329_2 , buf_splittern88ton117N329_N329_1 , buf_splitterfromn90_n125_3 , buf_splitterfromn90_n125_2 , buf_splitterfromn90_n125_1 , buf_splitterfromn93_n141_3 , buf_splitterfromn93_n141_2 , buf_splitterfromn93_n141_1 , buf_splitterfromn96_n127_3 , buf_splitterfromn96_n127_2 , buf_splitterfromn96_n127_1 , buf_splitterfromn101_n148_4 , buf_splitterfromn101_n148_3 , buf_splitterfromn101_n148_2 , buf_splitterfromn101_n148_1 , buf_splitterfromn104_n136_3 , buf_splitterfromn104_n136_2 , buf_splitterfromn104_n136_1 , buf_splitterfromn108_n138_4 , buf_splitterfromn108_n138_3 , buf_splitterfromn108_n138_2 , buf_splitterfromn108_n138_1 , buf_splitterfromn111_n131_4 , buf_splitterfromn111_n131_3 , buf_splitterfromn111_n131_2 , buf_splitterfromn111_n131_1 , buf_splitterfromn112_n132_3 , buf_splitterfromn112_n132_2 , buf_splitterfromn112_n132_1 , buf_splitterfromn115_n130_4 , buf_splitterfromn115_n130_3 , buf_splitterfromn115_n130_2 , buf_splitterfromn115_n130_1 , buf_splitterfromn118_n143_4 , buf_splitterfromn118_n143_3 , buf_splitterfromn118_n143_2 , buf_splitterfromn118_n143_1 , buf_splittern123ton140N370_N370_4 , buf_splittern123ton140N370_N370_3 , buf_splittern123ton140N370_N370_2 , buf_splittern123ton140N370_N370_1 , buf_splitterfromn125_n156_2 , buf_splitterfromn125_n156_1 , buf_splitterfromn127_n157_2 , buf_splitterfromn127_n157_1 , buf_splitterfromn134_N430_1 , buf_splitterfromn138_n152_1 , splitterfromN1 , splitterfromN102 , splitterfromN105 , splitterfromN108 , splitterfromN11 , splitterfromN112 , splitterfromN115 , splitterfromN14 , splitterfromN17 , splitterfromN21 , splitterfromN27 , splitterfromN30 , splitterfromN34 , splitterfromN37 , splitterfromN4 , splitterfromN40 , splitterfromN43 , splitterfromN47 , splitterfromN50 , splitterfromN53 , splitterfromN56 , splitterfromN60 , splitterfromN69 , splitterfromN73 , splitterfromN76 , splitterfromN79 , splitterfromN8 , splitterfromN82 , splitterfromN86 , splitterfromN89 , splitterfromN92 , splitterfromN95 , splitterfromN99 , splitterfromn37 , splitterfromn45 , splittern53ton79N223 , splittern53ton54n64 , splittern53ton69N223 , splitterfromn55 , splitterfromn58 , splitterfromn62 , splitterfromn65 , splitterfromn70 , splitterfromn73 , splitterfromn77 , splitterfromn80 , splitterfromn83 , splittern88ton110N329 , splittern88ton100n114 , splittern88ton117N329 , splitterfromn90 , splitterfromn93 , splitterfromn96 , splitterfromn101 , splitterfromn104 , splitterfromn108 , splitterfromn111 , splitterfromn112 , splitterfromn115 , splitterfromn118 , splittern123ton124N370 , splittern123ton129n137 , splittern123ton140N370 , splitterfromn125 , splitterfromn127 , splitterfromn128 , splitterfromn130 , splittern133ton134n152 , splitterfromn134 , splitterfromn136 , splitterfromn138 , splitterfromn139 , splitterfromn141 ;

PI_AQFP N1_( clk_1 , N1 );
PI_AQFP N102_( clk_1 , N102 );
PI_AQFP N105_( clk_1 , N105 );
PI_AQFP N108_( clk_1 , N108 );
PI_AQFP N11_( clk_1 , N11 );
PI_AQFP N112_( clk_1 , N112 );
PI_AQFP N115_( clk_1 , N115 );
PI_AQFP N14_( clk_1 , N14 );
PI_AQFP N17_( clk_1 , N17 );
PI_AQFP N21_( clk_1 , N21 );
PI_AQFP N24_( clk_1 , N24 );
PI_AQFP N27_( clk_1 , N27 );
PI_AQFP N30_( clk_1 , N30 );
PI_AQFP N34_( clk_1 , N34 );
PI_AQFP N37_( clk_1 , N37 );
PI_AQFP N4_( clk_1 , N4 );
PI_AQFP N40_( clk_1 , N40 );
PI_AQFP N43_( clk_1 , N43 );
PI_AQFP N47_( clk_1 , N47 );
PI_AQFP N50_( clk_1 , N50 );
PI_AQFP N53_( clk_1 , N53 );
PI_AQFP N56_( clk_1 , N56 );
PI_AQFP N60_( clk_1 , N60 );
PI_AQFP N63_( clk_1 , N63 );
PI_AQFP N66_( clk_1 , N66 );
PI_AQFP N69_( clk_1 , N69 );
PI_AQFP N73_( clk_1 , N73 );
PI_AQFP N76_( clk_1 , N76 );
PI_AQFP N79_( clk_1 , N79 );
PI_AQFP N8_( clk_1 , N8 );
PI_AQFP N82_( clk_1 , N82 );
PI_AQFP N86_( clk_1 , N86 );
PI_AQFP N89_( clk_1 , N89 );
PI_AQFP N92_( clk_1 , N92 );
PI_AQFP N95_( clk_1 , N95 );
PI_AQFP N99_( clk_1 , N99 );
and_AQFP n37_( clk_4 , buf_N24_n37_1 , splitterfromN30 , 1 , 0 , n37 );
and_AQFP n38_( clk_6 , splitterfromN102 , splitterfromN108 , 1 , 0 , n38 );
or_AQFP n39_( clk_7 , splitterfromn37 , n38 , 0 , 0 , n39 );
and_AQFP n40_( clk_5 , splitterfromN1 , splitterfromN4 , 1 , 0 , n40 );
and_AQFP n41_( clk_4 , splitterfromN89 , splitterfromN95 , 1 , 0 , n41 );
and_AQFP n42_( clk_4 , splitterfromN76 , splitterfromN82 , 1 , 0 , n42 );
or_AQFP n43_( clk_5 , n41 , n42 , 0 , 0 , n43 );
or_AQFP n44_( clk_6 , n40 , n43 , 0 , 0 , n44 );
and_AQFP n45_( clk_3 , N63 , splitterfromN69 , 1 , 0 , n45 );
and_AQFP n46_( clk_4 , splitterfromN37 , splitterfromN43 , 1 , 0 , n46 );
or_AQFP n47_( clk_5 , splitterfromn45 , n46 , 0 , 0 , n47 );
and_AQFP n48_( clk_4 , splitterfromN50 , splitterfromN56 , 1 , 0 , n48 );
and_AQFP n49_( clk_4 , splitterfromN11 , splitterfromN17 , 1 , 0 , n49 );
or_AQFP n50_( clk_5 , n48 , n49 , 0 , 0 , n50 );
or_AQFP n51_( clk_6 , n47 , n50 , 0 , 0 , n51 );
or_AQFP n52_( clk_7 , n44 , n51 , 0 , 0 , n52 );
or_AQFP n53_( clk_8 , n39 , n52 , 0 , 0 , n53 );
and_AQFP n54_( clk_3 , buf_splitterfromN102_n54_1 , splittern53ton54n64 , 0 , 0 , n54 );
and_AQFP n55_( clk_4 , buf_splitterfromN108_n55_1 , n54 , 0 , 1 , n55 );
and_AQFP n56_( clk_6 , splitterfromN112 , splitterfromn55 , 1 , 0 , n56 );
and_AQFP n57_( clk_3 , buf_splitterfromN76_n57_1 , splittern53ton54n64 , 0 , 0 , n57 );
and_AQFP n58_( clk_4 , buf_splitterfromN82_n58_1 , n57 , 0 , 1 , n58 );
and_AQFP n59_( clk_6 , splitterfromN86 , splitterfromn58 , 1 , 0 , n59 );
or_AQFP n60_( clk_7 , n56 , n59 , 0 , 0 , n60 );
and_AQFP n61_( clk_3 , buf_splitterfromN30_n61_1 , splittern53ton54n64 , 0 , 1 , n61 );
or_AQFP n62_( clk_4 , buf_splitterfromn37_n62_1 , n61 , 0 , 0 , n62 );
and_AQFP n63_( clk_6 , splitterfromN34 , splitterfromn62 , 1 , 0 , n63 );
and_AQFP n64_( clk_3 , buf_splitterfromN11_n64_1 , splittern53ton54n64 , 0 , 0 , n64 );
and_AQFP n65_( clk_4 , buf_splitterfromN17_n65_1 , n64 , 0 , 1 , n65 );
and_AQFP n66_( clk_6 , splitterfromN21 , splitterfromn65 , 1 , 0 , n66 );
or_AQFP n67_( clk_7 , n63 , n66 , 0 , 0 , n67 );
or_AQFP n68_( clk_8 , n60 , n67 , 0 , 0 , n68 );
and_AQFP n69_( clk_3 , buf_splitterfromN1_n69_1 , splittern53ton69N223 , 0 , 0 , n69 );
and_AQFP n70_( clk_4 , buf_splitterfromN4_n70_1 , n69 , 0 , 1 , n70 );
and_AQFP n71_( clk_6 , splitterfromN8 , splitterfromn70 , 1 , 0 , n71 );
and_AQFP n72_( clk_3 , buf_splitterfromN89_n72_1 , splittern53ton69N223 , 0 , 0 , n72 );
and_AQFP n73_( clk_4 , buf_splitterfromN95_n73_1 , n72 , 0 , 1 , n73 );
and_AQFP n74_( clk_6 , splitterfromN99 , splitterfromn73 , 1 , 0 , n74 );
or_AQFP n75_( clk_7 , n71 , n74 , 0 , 0 , n75 );
and_AQFP n76_( clk_3 , buf_splitterfromN50_n76_1 , splittern53ton69N223 , 0 , 0 , n76 );
and_AQFP n77_( clk_4 , buf_splitterfromN56_n77_1 , n76 , 0 , 1 , n77 );
and_AQFP n78_( clk_6 , splitterfromN60 , splitterfromn77 , 1 , 0 , n78 );
and_AQFP n79_( clk_2 , buf_splitterfromN69_n79_1 , splittern53ton79N223 , 0 , 1 , n79 );
or_AQFP n80_( clk_3 , buf_splitterfromn45_n80_1 , n79 , 0 , 0 , n80 );
and_AQFP n81_( clk_5 , splitterfromN73 , splitterfromn80 , 1 , 0 , n81 );
and_AQFP n82_( clk_2 , buf_splitterfromN37_n82_1 , splittern53ton79N223 , 0 , 0 , n82 );
and_AQFP n83_( clk_3 , buf_splitterfromN43_n83_1 , n82 , 0 , 1 , n83 );
and_AQFP n84_( clk_5 , splitterfromN47 , splitterfromn83 , 1 , 0 , n84 );
or_AQFP n85_( clk_6 , n81 , n84 , 0 , 0 , n85 );
or_AQFP n86_( clk_7 , n78 , n85 , 0 , 0 , n86 );
or_AQFP n87_( clk_8 , n75 , n86 , 0 , 0 , n87 );
or_AQFP n88_( clk_1 , n68 , n87 , 0 , 0 , n88 );
and_AQFP n89_( clk_4 , buf_splitterfromN34_n89_1 , splittern88ton117N329 , 0 , 0 , n89 );
and_AQFP n90_( clk_5 , buf_splitterfromn62_n90_1 , n89 , 0 , 1 , n90 );
and_AQFP n91_( clk_8 , splitterfromN40 , splitterfromn90 , 1 , 0 , n91 );
and_AQFP n92_( clk_3 , buf_splitterfromN99_n92_1 , splittern88ton110N329 , 0 , 0 , n92 );
and_AQFP n93_( clk_5 , buf_splitterfromn73_n93_1 , n92 , 0 , 1 , n93 );
and_AQFP n94_( clk_8 , splitterfromN105 , splitterfromn93 , 1 , 0 , n94 );
and_AQFP n95_( clk_4 , buf_splitterfromN21_n95_1 , splittern88ton117N329 , 0 , 0 , n95 );
and_AQFP n96_( clk_5 , buf_splitterfromn65_n96_1 , n95 , 0 , 1 , n96 );
and_AQFP n97_( clk_8 , splitterfromN27 , splitterfromn96 , 1 , 0 , n97 );
or_AQFP n98_( clk_1 , n94 , n97 , 0 , 0 , n98 );
or_AQFP n99_( clk_2 , n91 , n98 , 0 , 0 , n99 );
and_AQFP n100_( clk_4 , buf_splitterfromN8_n100_1 , splittern88ton100n114 , 0 , 0 , n100 );
and_AQFP n101_( clk_5 , buf_splitterfromn70_n101_1 , n100 , 0 , 1 , n101 );
and_AQFP n102_( clk_8 , splitterfromN14 , splitterfromn101 , 1 , 0 , n102 );
and_AQFP n103_( clk_4 , buf_splitterfromN86_n103_1 , splittern88ton100n114 , 0 , 0 , n103 );
and_AQFP n104_( clk_5 , buf_splitterfromn58_n104_1 , n103 , 0 , 1 , n104 );
and_AQFP n105_( clk_8 , splitterfromN92 , splitterfromn104 , 1 , 0 , n105 );
or_AQFP n106_( clk_1 , n102 , n105 , 0 , 0 , n106 );
and_AQFP n107_( clk_4 , buf_splitterfromN73_n107_1 , splittern88ton100n114 , 0 , 0 , n107 );
and_AQFP n108_( clk_5 , buf_splitterfromn80_n108_1 , n107 , 0 , 1 , n108 );
and_AQFP n109_( clk_7 , splitterfromN79 , splitterfromn108 , 1 , 0 , n109 );
and_AQFP n110_( clk_3 , buf_splitterfromN60_n110_1 , splittern88ton110N329 , 0 , 0 , n110 );
and_AQFP n111_( clk_4 , buf_splitterfromn77_n111_1 , n110 , 0 , 1 , n111 );
and_AQFP n112_( clk_6 , buf_N66_n112_1 , splitterfromn111 , 1 , 0 , n112 );
or_AQFP n113_( clk_8 , n109 , splitterfromn112 , 0 , 0 , n113 );
and_AQFP n114_( clk_4 , buf_splitterfromN47_n114_1 , splittern88ton100n114 , 0 , 0 , n114 );
and_AQFP n115_( clk_5 , buf_splitterfromn83_n115_1 , n114 , 0 , 1 , n115 );
and_AQFP n116_( clk_7 , splitterfromN53 , splitterfromn115 , 1 , 0 , n116 );
and_AQFP n117_( clk_4 , buf_splitterfromN112_n117_1 , splittern88ton117N329 , 0 , 0 , n117 );
and_AQFP n118_( clk_5 , buf_splitterfromn55_n118_1 , n117 , 0 , 1 , n118 );
and_AQFP n119_( clk_7 , splitterfromN115 , splitterfromn118 , 1 , 0 , n119 );
or_AQFP n120_( clk_8 , n116 , n119 , 0 , 0 , n120 );
or_AQFP n121_( clk_1 , n113 , n120 , 0 , 0 , n121 );
or_AQFP n122_( clk_2 , n106 , n121 , 0 , 0 , n122 );
or_AQFP n123_( clk_3 , n99 , n122 , 0 , 0 , n123 );
and_AQFP n124_( clk_5 , buf_splitterfromN40_n124_1 , splittern123ton124N370 , 0 , 0 , n124 );
and_AQFP n125_( clk_6 , buf_splitterfromn90_n125_1 , n124 , 0 , 1 , n125 );
and_AQFP n126_( clk_5 , buf_splitterfromN27_n126_1 , splittern123ton124N370 , 0 , 0 , n126 );
and_AQFP n127_( clk_6 , buf_splitterfromn96_n127_1 , n126 , 0 , 1 , n127 );
or_AQFP n128_( clk_1 , splitterfromn125 , splitterfromn127 , 0 , 0 , n128 );
and_AQFP n129_( clk_6 , buf_splitterfromN53_n129_1 , splittern123ton129n137 , 0 , 0 , n129 );
and_AQFP n130_( clk_7 , buf_splitterfromn115_n130_1 , n129 , 0 , 1 , n130 );
and_AQFP n131_( clk_6 , buf_splitterfromn111_n131_1 , splittern123ton129n137 , 0 , 1 , n131 );
or_AQFP n132_( clk_7 , buf_splitterfromn112_n132_1 , n131 , 0 , 0 , n132 );
or_AQFP n133_( clk_1 , splitterfromn130 , n132 , 0 , 0 , n133 );
or_AQFP n134_( clk_3 , splitterfromn128 , splittern133ton134n152 , 0 , 0 , n134 );
and_AQFP n135_( clk_6 , buf_splitterfromN92_n135_1 , splittern123ton129n137 , 0 , 0 , n135 );
and_AQFP n136_( clk_7 , buf_splitterfromn104_n136_1 , n135 , 0 , 1 , n136 );
and_AQFP n137_( clk_6 , buf_splitterfromN79_n137_1 , splittern123ton129n137 , 0 , 0 , n137 );
and_AQFP n138_( clk_7 , buf_splitterfromn108_n138_1 , n137 , 0 , 1 , n138 );
or_AQFP n139_( clk_1 , splitterfromn136 , splitterfromn138 , 0 , 0 , n139 );
and_AQFP n140_( clk_6 , buf_splitterfromN105_n140_1 , splittern123ton140N370 , 0 , 0 , n140 );
and_AQFP n141_( clk_7 , buf_splitterfromn93_n141_1 , n140 , 0 , 1 , n141 );
and_AQFP n142_( clk_6 , buf_splitterfromN115_n142_1 , splittern123ton140N370 , 0 , 0 , n142 );
and_AQFP n143_( clk_7 , buf_splitterfromn118_n143_1 , n142 , 0 , 1 , n143 );
or_AQFP n144_( clk_1 , splitterfromn141 , n143 , 0 , 0 , n144 );
or_AQFP n145_( clk_3 , splitterfromn139 , n144 , 0 , 0 , n145 );
or_AQFP n146_( clk_5 , splitterfromn134 , n145 , 0 , 0 , n146 );
and_AQFP n147_( clk_6 , buf_splitterfromN14_n147_1 , splittern123ton140N370 , 0 , 0 , n147 );
and_AQFP n148_( clk_8 , buf_splitterfromn101_n148_1 , n147 , 0 , 1 , n148 );
and_AQFP n149_( clk_6 , n146 , buf_n148_n149_1 , 0 , 1 , n149 );
and_AQFP n150_( clk_3 , splittern133ton134n152 , splitterfromn139 , 1 , 0 , n150 );
or_AQFP n151_( clk_4 , splitterfromn128 , n150 , 0 , 0 , n151 );
and_AQFP n152_( clk_3 , splittern133ton134n152 , buf_splitterfromn138_n152_1 , 1 , 0 , n152 );
and_AQFP n153_( clk_1 , splitterfromn136 , splitterfromn141 , 1 , 0 , n153 );
or_AQFP n154_( clk_2 , splitterfromn130 , n153 , 0 , 0 , n154 );
or_AQFP n155_( clk_4 , n152 , n154 , 0 , 0 , n155 );
and_AQFP n156_( clk_5 , buf_splitterfromn125_n156_1 , n155 , 1 , 0 , n156 );
or_AQFP n157_( clk_6 , buf_splitterfromn127_n157_1 , n156 , 0 , 0 , n157 );
PO_AQFP N223_( clk_7 , buf_splittern53ton69N223_N223_1 , 0 , N223 );
PO_AQFP N329_( clk_7 , buf_splittern88ton117N329_N329_1 , 0 , N329 );
PO_AQFP N370_( clk_7 , buf_splittern123ton140N370_N370_1 , 0 , N370 );
PO_AQFP N421_( clk_7 , n149 , 0 , N421 );
PO_AQFP N430_( clk_7 , buf_splitterfromn134_N430_1 , 0 , N430 );
PO_AQFP N431_( clk_7 , buf_n151_N431_1 , 0 , N431 );
PO_AQFP N432_( clk_7 , n157 , 0 , N432 );
buf_AQFP buf_N102_splitterfromN102_1_( clk_3 , N102 , 0 , buf_N102_splitterfromN102_1 );
buf_AQFP buf_N105_splitterfromN105_10_( clk_3 , N105 , 0 , buf_N105_splitterfromN105_10 );
buf_AQFP buf_N105_splitterfromN105_9_( clk_5 , buf_N105_splitterfromN105_10 , 0 , buf_N105_splitterfromN105_9 );
buf_AQFP buf_N105_splitterfromN105_8_( clk_7 , buf_N105_splitterfromN105_9 , 0 , buf_N105_splitterfromN105_8 );
buf_AQFP buf_N105_splitterfromN105_7_( clk_1 , buf_N105_splitterfromN105_8 , 0 , buf_N105_splitterfromN105_7 );
buf_AQFP buf_N105_splitterfromN105_6_( clk_3 , buf_N105_splitterfromN105_7 , 0 , buf_N105_splitterfromN105_6 );
buf_AQFP buf_N105_splitterfromN105_5_( clk_5 , buf_N105_splitterfromN105_6 , 0 , buf_N105_splitterfromN105_5 );
buf_AQFP buf_N105_splitterfromN105_4_( clk_7 , buf_N105_splitterfromN105_5 , 0 , buf_N105_splitterfromN105_4 );
buf_AQFP buf_N105_splitterfromN105_3_( clk_1 , buf_N105_splitterfromN105_4 , 0 , buf_N105_splitterfromN105_3 );
buf_AQFP buf_N105_splitterfromN105_2_( clk_3 , buf_N105_splitterfromN105_3 , 0 , buf_N105_splitterfromN105_2 );
buf_AQFP buf_N105_splitterfromN105_1_( clk_5 , buf_N105_splitterfromN105_2 , 0 , buf_N105_splitterfromN105_1 );
buf_AQFP buf_N108_splitterfromN108_1_( clk_3 , N108 , 0 , buf_N108_splitterfromN108_1 );
buf_AQFP buf_N112_splitterfromN112_5_( clk_3 , N112 , 0 , buf_N112_splitterfromN112_5 );
buf_AQFP buf_N112_splitterfromN112_4_( clk_5 , buf_N112_splitterfromN112_5 , 0 , buf_N112_splitterfromN112_4 );
buf_AQFP buf_N112_splitterfromN112_3_( clk_7 , buf_N112_splitterfromN112_4 , 0 , buf_N112_splitterfromN112_3 );
buf_AQFP buf_N112_splitterfromN112_2_( clk_1 , buf_N112_splitterfromN112_3 , 0 , buf_N112_splitterfromN112_2 );
buf_AQFP buf_N112_splitterfromN112_1_( clk_3 , buf_N112_splitterfromN112_2 , 0 , buf_N112_splitterfromN112_1 );
buf_AQFP buf_N115_splitterfromN115_10_( clk_3 , N115 , 0 , buf_N115_splitterfromN115_10 );
buf_AQFP buf_N115_splitterfromN115_9_( clk_5 , buf_N115_splitterfromN115_10 , 0 , buf_N115_splitterfromN115_9 );
buf_AQFP buf_N115_splitterfromN115_8_( clk_7 , buf_N115_splitterfromN115_9 , 0 , buf_N115_splitterfromN115_8 );
buf_AQFP buf_N115_splitterfromN115_7_( clk_1 , buf_N115_splitterfromN115_8 , 0 , buf_N115_splitterfromN115_7 );
buf_AQFP buf_N115_splitterfromN115_6_( clk_3 , buf_N115_splitterfromN115_7 , 0 , buf_N115_splitterfromN115_6 );
buf_AQFP buf_N115_splitterfromN115_5_( clk_5 , buf_N115_splitterfromN115_6 , 0 , buf_N115_splitterfromN115_5 );
buf_AQFP buf_N115_splitterfromN115_4_( clk_7 , buf_N115_splitterfromN115_5 , 0 , buf_N115_splitterfromN115_4 );
buf_AQFP buf_N115_splitterfromN115_3_( clk_1 , buf_N115_splitterfromN115_4 , 0 , buf_N115_splitterfromN115_3 );
buf_AQFP buf_N115_splitterfromN115_2_( clk_3 , buf_N115_splitterfromN115_3 , 0 , buf_N115_splitterfromN115_2 );
buf_AQFP buf_N115_splitterfromN115_1_( clk_5 , buf_N115_splitterfromN115_2 , 0 , buf_N115_splitterfromN115_1 );
buf_AQFP buf_N14_splitterfromN14_10_( clk_3 , N14 , 0 , buf_N14_splitterfromN14_10 );
buf_AQFP buf_N14_splitterfromN14_9_( clk_5 , buf_N14_splitterfromN14_10 , 0 , buf_N14_splitterfromN14_9 );
buf_AQFP buf_N14_splitterfromN14_8_( clk_7 , buf_N14_splitterfromN14_9 , 0 , buf_N14_splitterfromN14_8 );
buf_AQFP buf_N14_splitterfromN14_7_( clk_1 , buf_N14_splitterfromN14_8 , 0 , buf_N14_splitterfromN14_7 );
buf_AQFP buf_N14_splitterfromN14_6_( clk_3 , buf_N14_splitterfromN14_7 , 0 , buf_N14_splitterfromN14_6 );
buf_AQFP buf_N14_splitterfromN14_5_( clk_5 , buf_N14_splitterfromN14_6 , 0 , buf_N14_splitterfromN14_5 );
buf_AQFP buf_N14_splitterfromN14_4_( clk_7 , buf_N14_splitterfromN14_5 , 0 , buf_N14_splitterfromN14_4 );
buf_AQFP buf_N14_splitterfromN14_3_( clk_1 , buf_N14_splitterfromN14_4 , 0 , buf_N14_splitterfromN14_3 );
buf_AQFP buf_N14_splitterfromN14_2_( clk_3 , buf_N14_splitterfromN14_3 , 0 , buf_N14_splitterfromN14_2 );
buf_AQFP buf_N14_splitterfromN14_1_( clk_5 , buf_N14_splitterfromN14_2 , 0 , buf_N14_splitterfromN14_1 );
buf_AQFP buf_N21_splitterfromN21_5_( clk_3 , N21 , 0 , buf_N21_splitterfromN21_5 );
buf_AQFP buf_N21_splitterfromN21_4_( clk_5 , buf_N21_splitterfromN21_5 , 0 , buf_N21_splitterfromN21_4 );
buf_AQFP buf_N21_splitterfromN21_3_( clk_7 , buf_N21_splitterfromN21_4 , 0 , buf_N21_splitterfromN21_3 );
buf_AQFP buf_N21_splitterfromN21_2_( clk_1 , buf_N21_splitterfromN21_3 , 0 , buf_N21_splitterfromN21_2 );
buf_AQFP buf_N21_splitterfromN21_1_( clk_3 , buf_N21_splitterfromN21_2 , 0 , buf_N21_splitterfromN21_1 );
buf_AQFP buf_N24_n37_1_( clk_3 , N24 , 0 , buf_N24_n37_1 );
buf_AQFP buf_N27_splitterfromN27_10_( clk_3 , N27 , 0 , buf_N27_splitterfromN27_10 );
buf_AQFP buf_N27_splitterfromN27_9_( clk_5 , buf_N27_splitterfromN27_10 , 0 , buf_N27_splitterfromN27_9 );
buf_AQFP buf_N27_splitterfromN27_8_( clk_7 , buf_N27_splitterfromN27_9 , 0 , buf_N27_splitterfromN27_8 );
buf_AQFP buf_N27_splitterfromN27_7_( clk_1 , buf_N27_splitterfromN27_8 , 0 , buf_N27_splitterfromN27_7 );
buf_AQFP buf_N27_splitterfromN27_6_( clk_3 , buf_N27_splitterfromN27_7 , 0 , buf_N27_splitterfromN27_6 );
buf_AQFP buf_N27_splitterfromN27_5_( clk_5 , buf_N27_splitterfromN27_6 , 0 , buf_N27_splitterfromN27_5 );
buf_AQFP buf_N27_splitterfromN27_4_( clk_7 , buf_N27_splitterfromN27_5 , 0 , buf_N27_splitterfromN27_4 );
buf_AQFP buf_N27_splitterfromN27_3_( clk_1 , buf_N27_splitterfromN27_4 , 0 , buf_N27_splitterfromN27_3 );
buf_AQFP buf_N27_splitterfromN27_2_( clk_3 , buf_N27_splitterfromN27_3 , 0 , buf_N27_splitterfromN27_2 );
buf_AQFP buf_N27_splitterfromN27_1_( clk_5 , buf_N27_splitterfromN27_2 , 0 , buf_N27_splitterfromN27_1 );
buf_AQFP buf_N34_splitterfromN34_5_( clk_3 , N34 , 0 , buf_N34_splitterfromN34_5 );
buf_AQFP buf_N34_splitterfromN34_4_( clk_5 , buf_N34_splitterfromN34_5 , 0 , buf_N34_splitterfromN34_4 );
buf_AQFP buf_N34_splitterfromN34_3_( clk_7 , buf_N34_splitterfromN34_4 , 0 , buf_N34_splitterfromN34_3 );
buf_AQFP buf_N34_splitterfromN34_2_( clk_1 , buf_N34_splitterfromN34_3 , 0 , buf_N34_splitterfromN34_2 );
buf_AQFP buf_N34_splitterfromN34_1_( clk_3 , buf_N34_splitterfromN34_2 , 0 , buf_N34_splitterfromN34_1 );
buf_AQFP buf_N4_splitterfromN4_1_( clk_3 , N4 , 0 , buf_N4_splitterfromN4_1 );
buf_AQFP buf_N40_splitterfromN40_10_( clk_3 , N40 , 0 , buf_N40_splitterfromN40_10 );
buf_AQFP buf_N40_splitterfromN40_9_( clk_5 , buf_N40_splitterfromN40_10 , 0 , buf_N40_splitterfromN40_9 );
buf_AQFP buf_N40_splitterfromN40_8_( clk_7 , buf_N40_splitterfromN40_9 , 0 , buf_N40_splitterfromN40_8 );
buf_AQFP buf_N40_splitterfromN40_7_( clk_1 , buf_N40_splitterfromN40_8 , 0 , buf_N40_splitterfromN40_7 );
buf_AQFP buf_N40_splitterfromN40_6_( clk_3 , buf_N40_splitterfromN40_7 , 0 , buf_N40_splitterfromN40_6 );
buf_AQFP buf_N40_splitterfromN40_5_( clk_5 , buf_N40_splitterfromN40_6 , 0 , buf_N40_splitterfromN40_5 );
buf_AQFP buf_N40_splitterfromN40_4_( clk_7 , buf_N40_splitterfromN40_5 , 0 , buf_N40_splitterfromN40_4 );
buf_AQFP buf_N40_splitterfromN40_3_( clk_1 , buf_N40_splitterfromN40_4 , 0 , buf_N40_splitterfromN40_3 );
buf_AQFP buf_N40_splitterfromN40_2_( clk_3 , buf_N40_splitterfromN40_3 , 0 , buf_N40_splitterfromN40_2 );
buf_AQFP buf_N40_splitterfromN40_1_( clk_5 , buf_N40_splitterfromN40_2 , 0 , buf_N40_splitterfromN40_1 );
buf_AQFP buf_N47_splitterfromN47_5_( clk_3 , N47 , 0 , buf_N47_splitterfromN47_5 );
buf_AQFP buf_N47_splitterfromN47_4_( clk_5 , buf_N47_splitterfromN47_5 , 0 , buf_N47_splitterfromN47_4 );
buf_AQFP buf_N47_splitterfromN47_3_( clk_7 , buf_N47_splitterfromN47_4 , 0 , buf_N47_splitterfromN47_3 );
buf_AQFP buf_N47_splitterfromN47_2_( clk_1 , buf_N47_splitterfromN47_3 , 0 , buf_N47_splitterfromN47_2 );
buf_AQFP buf_N47_splitterfromN47_1_( clk_3 , buf_N47_splitterfromN47_2 , 0 , buf_N47_splitterfromN47_1 );
buf_AQFP buf_N53_splitterfromN53_10_( clk_3 , N53 , 0 , buf_N53_splitterfromN53_10 );
buf_AQFP buf_N53_splitterfromN53_9_( clk_5 , buf_N53_splitterfromN53_10 , 0 , buf_N53_splitterfromN53_9 );
buf_AQFP buf_N53_splitterfromN53_8_( clk_7 , buf_N53_splitterfromN53_9 , 0 , buf_N53_splitterfromN53_8 );
buf_AQFP buf_N53_splitterfromN53_7_( clk_1 , buf_N53_splitterfromN53_8 , 0 , buf_N53_splitterfromN53_7 );
buf_AQFP buf_N53_splitterfromN53_6_( clk_3 , buf_N53_splitterfromN53_7 , 0 , buf_N53_splitterfromN53_6 );
buf_AQFP buf_N53_splitterfromN53_5_( clk_5 , buf_N53_splitterfromN53_6 , 0 , buf_N53_splitterfromN53_5 );
buf_AQFP buf_N53_splitterfromN53_4_( clk_7 , buf_N53_splitterfromN53_5 , 0 , buf_N53_splitterfromN53_4 );
buf_AQFP buf_N53_splitterfromN53_3_( clk_1 , buf_N53_splitterfromN53_4 , 0 , buf_N53_splitterfromN53_3 );
buf_AQFP buf_N53_splitterfromN53_2_( clk_3 , buf_N53_splitterfromN53_3 , 0 , buf_N53_splitterfromN53_2 );
buf_AQFP buf_N53_splitterfromN53_1_( clk_5 , buf_N53_splitterfromN53_2 , 0 , buf_N53_splitterfromN53_1 );
buf_AQFP buf_N60_splitterfromN60_5_( clk_3 , N60 , 0 , buf_N60_splitterfromN60_5 );
buf_AQFP buf_N60_splitterfromN60_4_( clk_5 , buf_N60_splitterfromN60_5 , 0 , buf_N60_splitterfromN60_4 );
buf_AQFP buf_N60_splitterfromN60_3_( clk_7 , buf_N60_splitterfromN60_4 , 0 , buf_N60_splitterfromN60_3 );
buf_AQFP buf_N60_splitterfromN60_2_( clk_1 , buf_N60_splitterfromN60_3 , 0 , buf_N60_splitterfromN60_2 );
buf_AQFP buf_N60_splitterfromN60_1_( clk_3 , buf_N60_splitterfromN60_2 , 0 , buf_N60_splitterfromN60_1 );
buf_AQFP buf_N66_n112_10_( clk_3 , N66 , 0 , buf_N66_n112_10 );
buf_AQFP buf_N66_n112_9_( clk_5 , buf_N66_n112_10 , 0 , buf_N66_n112_9 );
buf_AQFP buf_N66_n112_8_( clk_7 , buf_N66_n112_9 , 0 , buf_N66_n112_8 );
buf_AQFP buf_N66_n112_7_( clk_1 , buf_N66_n112_8 , 0 , buf_N66_n112_7 );
buf_AQFP buf_N66_n112_6_( clk_3 , buf_N66_n112_7 , 0 , buf_N66_n112_6 );
buf_AQFP buf_N66_n112_5_( clk_5 , buf_N66_n112_6 , 0 , buf_N66_n112_5 );
buf_AQFP buf_N66_n112_4_( clk_7 , buf_N66_n112_5 , 0 , buf_N66_n112_4 );
buf_AQFP buf_N66_n112_3_( clk_1 , buf_N66_n112_4 , 0 , buf_N66_n112_3 );
buf_AQFP buf_N66_n112_2_( clk_3 , buf_N66_n112_3 , 0 , buf_N66_n112_2 );
buf_AQFP buf_N66_n112_1_( clk_5 , buf_N66_n112_2 , 0 , buf_N66_n112_1 );
buf_AQFP buf_N73_splitterfromN73_5_( clk_3 , N73 , 0 , buf_N73_splitterfromN73_5 );
buf_AQFP buf_N73_splitterfromN73_4_( clk_5 , buf_N73_splitterfromN73_5 , 0 , buf_N73_splitterfromN73_4 );
buf_AQFP buf_N73_splitterfromN73_3_( clk_7 , buf_N73_splitterfromN73_4 , 0 , buf_N73_splitterfromN73_3 );
buf_AQFP buf_N73_splitterfromN73_2_( clk_1 , buf_N73_splitterfromN73_3 , 0 , buf_N73_splitterfromN73_2 );
buf_AQFP buf_N73_splitterfromN73_1_( clk_3 , buf_N73_splitterfromN73_2 , 0 , buf_N73_splitterfromN73_1 );
buf_AQFP buf_N79_splitterfromN79_10_( clk_3 , N79 , 0 , buf_N79_splitterfromN79_10 );
buf_AQFP buf_N79_splitterfromN79_9_( clk_5 , buf_N79_splitterfromN79_10 , 0 , buf_N79_splitterfromN79_9 );
buf_AQFP buf_N79_splitterfromN79_8_( clk_7 , buf_N79_splitterfromN79_9 , 0 , buf_N79_splitterfromN79_8 );
buf_AQFP buf_N79_splitterfromN79_7_( clk_1 , buf_N79_splitterfromN79_8 , 0 , buf_N79_splitterfromN79_7 );
buf_AQFP buf_N79_splitterfromN79_6_( clk_3 , buf_N79_splitterfromN79_7 , 0 , buf_N79_splitterfromN79_6 );
buf_AQFP buf_N79_splitterfromN79_5_( clk_5 , buf_N79_splitterfromN79_6 , 0 , buf_N79_splitterfromN79_5 );
buf_AQFP buf_N79_splitterfromN79_4_( clk_7 , buf_N79_splitterfromN79_5 , 0 , buf_N79_splitterfromN79_4 );
buf_AQFP buf_N79_splitterfromN79_3_( clk_1 , buf_N79_splitterfromN79_4 , 0 , buf_N79_splitterfromN79_3 );
buf_AQFP buf_N79_splitterfromN79_2_( clk_3 , buf_N79_splitterfromN79_3 , 0 , buf_N79_splitterfromN79_2 );
buf_AQFP buf_N79_splitterfromN79_1_( clk_5 , buf_N79_splitterfromN79_2 , 0 , buf_N79_splitterfromN79_1 );
buf_AQFP buf_N8_splitterfromN8_5_( clk_3 , N8 , 0 , buf_N8_splitterfromN8_5 );
buf_AQFP buf_N8_splitterfromN8_4_( clk_5 , buf_N8_splitterfromN8_5 , 0 , buf_N8_splitterfromN8_4 );
buf_AQFP buf_N8_splitterfromN8_3_( clk_7 , buf_N8_splitterfromN8_4 , 0 , buf_N8_splitterfromN8_3 );
buf_AQFP buf_N8_splitterfromN8_2_( clk_1 , buf_N8_splitterfromN8_3 , 0 , buf_N8_splitterfromN8_2 );
buf_AQFP buf_N8_splitterfromN8_1_( clk_3 , buf_N8_splitterfromN8_2 , 0 , buf_N8_splitterfromN8_1 );
buf_AQFP buf_N86_splitterfromN86_5_( clk_3 , N86 , 0 , buf_N86_splitterfromN86_5 );
buf_AQFP buf_N86_splitterfromN86_4_( clk_5 , buf_N86_splitterfromN86_5 , 0 , buf_N86_splitterfromN86_4 );
buf_AQFP buf_N86_splitterfromN86_3_( clk_7 , buf_N86_splitterfromN86_4 , 0 , buf_N86_splitterfromN86_3 );
buf_AQFP buf_N86_splitterfromN86_2_( clk_1 , buf_N86_splitterfromN86_3 , 0 , buf_N86_splitterfromN86_2 );
buf_AQFP buf_N86_splitterfromN86_1_( clk_3 , buf_N86_splitterfromN86_2 , 0 , buf_N86_splitterfromN86_1 );
buf_AQFP buf_N92_splitterfromN92_10_( clk_3 , N92 , 0 , buf_N92_splitterfromN92_10 );
buf_AQFP buf_N92_splitterfromN92_9_( clk_5 , buf_N92_splitterfromN92_10 , 0 , buf_N92_splitterfromN92_9 );
buf_AQFP buf_N92_splitterfromN92_8_( clk_7 , buf_N92_splitterfromN92_9 , 0 , buf_N92_splitterfromN92_8 );
buf_AQFP buf_N92_splitterfromN92_7_( clk_1 , buf_N92_splitterfromN92_8 , 0 , buf_N92_splitterfromN92_7 );
buf_AQFP buf_N92_splitterfromN92_6_( clk_3 , buf_N92_splitterfromN92_7 , 0 , buf_N92_splitterfromN92_6 );
buf_AQFP buf_N92_splitterfromN92_5_( clk_5 , buf_N92_splitterfromN92_6 , 0 , buf_N92_splitterfromN92_5 );
buf_AQFP buf_N92_splitterfromN92_4_( clk_7 , buf_N92_splitterfromN92_5 , 0 , buf_N92_splitterfromN92_4 );
buf_AQFP buf_N92_splitterfromN92_3_( clk_1 , buf_N92_splitterfromN92_4 , 0 , buf_N92_splitterfromN92_3 );
buf_AQFP buf_N92_splitterfromN92_2_( clk_3 , buf_N92_splitterfromN92_3 , 0 , buf_N92_splitterfromN92_2 );
buf_AQFP buf_N92_splitterfromN92_1_( clk_5 , buf_N92_splitterfromN92_2 , 0 , buf_N92_splitterfromN92_1 );
buf_AQFP buf_N99_splitterfromN99_5_( clk_3 , N99 , 0 , buf_N99_splitterfromN99_5 );
buf_AQFP buf_N99_splitterfromN99_4_( clk_5 , buf_N99_splitterfromN99_5 , 0 , buf_N99_splitterfromN99_4 );
buf_AQFP buf_N99_splitterfromN99_3_( clk_7 , buf_N99_splitterfromN99_4 , 0 , buf_N99_splitterfromN99_3 );
buf_AQFP buf_N99_splitterfromN99_2_( clk_1 , buf_N99_splitterfromN99_3 , 0 , buf_N99_splitterfromN99_2 );
buf_AQFP buf_N99_splitterfromN99_1_( clk_3 , buf_N99_splitterfromN99_2 , 0 , buf_N99_splitterfromN99_1 );
buf_AQFP buf_n148_n149_2_( clk_2 , n148 , 0 , buf_n148_n149_2 );
buf_AQFP buf_n148_n149_1_( clk_4 , buf_n148_n149_2 , 0 , buf_n148_n149_1 );
buf_AQFP buf_n151_N431_1_( clk_6 , n151 , 0 , buf_n151_N431_1 );
buf_AQFP buf_splitterfromN1_n69_3_( clk_5 , splitterfromN1 , 0 , buf_splitterfromN1_n69_3 );
buf_AQFP buf_splitterfromN1_n69_2_( clk_7 , buf_splitterfromN1_n69_3 , 0 , buf_splitterfromN1_n69_2 );
buf_AQFP buf_splitterfromN1_n69_1_( clk_1 , buf_splitterfromN1_n69_2 , 0 , buf_splitterfromN1_n69_1 );
buf_AQFP buf_splitterfromN102_n54_2_( clk_7 , splitterfromN102 , 0 , buf_splitterfromN102_n54_2 );
buf_AQFP buf_splitterfromN102_n54_1_( clk_1 , buf_splitterfromN102_n54_2 , 0 , buf_splitterfromN102_n54_1 );
buf_AQFP buf_splitterfromN105_n140_3_( clk_1 , splitterfromN105 , 0 , buf_splitterfromN105_n140_3 );
buf_AQFP buf_splitterfromN105_n140_2_( clk_3 , buf_splitterfromN105_n140_3 , 0 , buf_splitterfromN105_n140_2 );
buf_AQFP buf_splitterfromN105_n140_1_( clk_5 , buf_splitterfromN105_n140_2 , 0 , buf_splitterfromN105_n140_1 );
buf_AQFP buf_splitterfromN108_n55_3_( clk_7 , splitterfromN108 , 0 , buf_splitterfromN108_n55_3 );
buf_AQFP buf_splitterfromN108_n55_2_( clk_1 , buf_splitterfromN108_n55_3 , 0 , buf_splitterfromN108_n55_2 );
buf_AQFP buf_splitterfromN108_n55_1_( clk_3 , buf_splitterfromN108_n55_2 , 0 , buf_splitterfromN108_n55_1 );
buf_AQFP buf_splitterfromN11_n64_3_( clk_5 , splitterfromN11 , 0 , buf_splitterfromN11_n64_3 );
buf_AQFP buf_splitterfromN11_n64_2_( clk_7 , buf_splitterfromN11_n64_3 , 0 , buf_splitterfromN11_n64_2 );
buf_AQFP buf_splitterfromN11_n64_1_( clk_1 , buf_splitterfromN11_n64_2 , 0 , buf_splitterfromN11_n64_1 );
buf_AQFP buf_splitterfromN112_n117_3_( clk_6 , splitterfromN112 , 0 , buf_splitterfromN112_n117_3 );
buf_AQFP buf_splitterfromN112_n117_2_( clk_8 , buf_splitterfromN112_n117_3 , 0 , buf_splitterfromN112_n117_2 );
buf_AQFP buf_splitterfromN112_n117_1_( clk_2 , buf_splitterfromN112_n117_2 , 0 , buf_splitterfromN112_n117_1 );
buf_AQFP buf_splitterfromN115_n142_3_( clk_8 , splitterfromN115 , 0 , buf_splitterfromN115_n142_3 );
buf_AQFP buf_splitterfromN115_n142_2_( clk_2 , buf_splitterfromN115_n142_3 , 0 , buf_splitterfromN115_n142_2 );
buf_AQFP buf_splitterfromN115_n142_1_( clk_4 , buf_splitterfromN115_n142_2 , 0 , buf_splitterfromN115_n142_1 );
buf_AQFP buf_splitterfromN14_n147_3_( clk_1 , splitterfromN14 , 0 , buf_splitterfromN14_n147_3 );
buf_AQFP buf_splitterfromN14_n147_2_( clk_3 , buf_splitterfromN14_n147_3 , 0 , buf_splitterfromN14_n147_2 );
buf_AQFP buf_splitterfromN14_n147_1_( clk_5 , buf_splitterfromN14_n147_2 , 0 , buf_splitterfromN14_n147_1 );
buf_AQFP buf_splitterfromN17_n65_4_( clk_5 , splitterfromN17 , 0 , buf_splitterfromN17_n65_4 );
buf_AQFP buf_splitterfromN17_n65_3_( clk_7 , buf_splitterfromN17_n65_4 , 0 , buf_splitterfromN17_n65_3 );
buf_AQFP buf_splitterfromN17_n65_2_( clk_1 , buf_splitterfromN17_n65_3 , 0 , buf_splitterfromN17_n65_2 );
buf_AQFP buf_splitterfromN17_n65_1_( clk_3 , buf_splitterfromN17_n65_2 , 0 , buf_splitterfromN17_n65_1 );
buf_AQFP buf_splitterfromN21_n95_3_( clk_7 , splitterfromN21 , 0 , buf_splitterfromN21_n95_3 );
buf_AQFP buf_splitterfromN21_n95_2_( clk_1 , buf_splitterfromN21_n95_3 , 0 , buf_splitterfromN21_n95_2 );
buf_AQFP buf_splitterfromN21_n95_1_( clk_3 , buf_splitterfromN21_n95_2 , 0 , buf_splitterfromN21_n95_1 );
buf_AQFP buf_splitterfromN27_n126_2_( clk_1 , splitterfromN27 , 0 , buf_splitterfromN27_n126_2 );
buf_AQFP buf_splitterfromN27_n126_1_( clk_3 , buf_splitterfromN27_n126_2 , 0 , buf_splitterfromN27_n126_1 );
buf_AQFP buf_splitterfromN30_n61_3_( clk_5 , splitterfromN30 , 0 , buf_splitterfromN30_n61_3 );
buf_AQFP buf_splitterfromN30_n61_2_( clk_7 , buf_splitterfromN30_n61_3 , 0 , buf_splitterfromN30_n61_2 );
buf_AQFP buf_splitterfromN30_n61_1_( clk_1 , buf_splitterfromN30_n61_2 , 0 , buf_splitterfromN30_n61_1 );
buf_AQFP buf_splitterfromN34_n89_3_( clk_7 , splitterfromN34 , 0 , buf_splitterfromN34_n89_3 );
buf_AQFP buf_splitterfromN34_n89_2_( clk_1 , buf_splitterfromN34_n89_3 , 0 , buf_splitterfromN34_n89_2 );
buf_AQFP buf_splitterfromN34_n89_1_( clk_3 , buf_splitterfromN34_n89_2 , 0 , buf_splitterfromN34_n89_1 );
buf_AQFP buf_splitterfromN37_n82_3_( clk_5 , splitterfromN37 , 0 , buf_splitterfromN37_n82_3 );
buf_AQFP buf_splitterfromN37_n82_2_( clk_7 , buf_splitterfromN37_n82_3 , 0 , buf_splitterfromN37_n82_2 );
buf_AQFP buf_splitterfromN37_n82_1_( clk_1 , buf_splitterfromN37_n82_2 , 0 , buf_splitterfromN37_n82_1 );
buf_AQFP buf_splitterfromN4_n70_3_( clk_6 , splitterfromN4 , 0 , buf_splitterfromN4_n70_3 );
buf_AQFP buf_splitterfromN4_n70_2_( clk_8 , buf_splitterfromN4_n70_3 , 0 , buf_splitterfromN4_n70_2 );
buf_AQFP buf_splitterfromN4_n70_1_( clk_2 , buf_splitterfromN4_n70_2 , 0 , buf_splitterfromN4_n70_1 );
buf_AQFP buf_splitterfromN40_n124_2_( clk_1 , splitterfromN40 , 0 , buf_splitterfromN40_n124_2 );
buf_AQFP buf_splitterfromN40_n124_1_( clk_3 , buf_splitterfromN40_n124_2 , 0 , buf_splitterfromN40_n124_1 );
buf_AQFP buf_splitterfromN43_n83_3_( clk_5 , splitterfromN43 , 0 , buf_splitterfromN43_n83_3 );
buf_AQFP buf_splitterfromN43_n83_2_( clk_7 , buf_splitterfromN43_n83_3 , 0 , buf_splitterfromN43_n83_2 );
buf_AQFP buf_splitterfromN43_n83_1_( clk_1 , buf_splitterfromN43_n83_2 , 0 , buf_splitterfromN43_n83_1 );
buf_AQFP buf_splitterfromN47_n114_3_( clk_6 , splitterfromN47 , 0 , buf_splitterfromN47_n114_3 );
buf_AQFP buf_splitterfromN47_n114_2_( clk_8 , buf_splitterfromN47_n114_3 , 0 , buf_splitterfromN47_n114_2 );
buf_AQFP buf_splitterfromN47_n114_1_( clk_2 , buf_splitterfromN47_n114_2 , 0 , buf_splitterfromN47_n114_1 );
buf_AQFP buf_splitterfromN50_n76_3_( clk_5 , splitterfromN50 , 0 , buf_splitterfromN50_n76_3 );
buf_AQFP buf_splitterfromN50_n76_2_( clk_7 , buf_splitterfromN50_n76_3 , 0 , buf_splitterfromN50_n76_2 );
buf_AQFP buf_splitterfromN50_n76_1_( clk_1 , buf_splitterfromN50_n76_2 , 0 , buf_splitterfromN50_n76_1 );
buf_AQFP buf_splitterfromN53_n129_3_( clk_8 , splitterfromN53 , 0 , buf_splitterfromN53_n129_3 );
buf_AQFP buf_splitterfromN53_n129_2_( clk_2 , buf_splitterfromN53_n129_3 , 0 , buf_splitterfromN53_n129_2 );
buf_AQFP buf_splitterfromN53_n129_1_( clk_4 , buf_splitterfromN53_n129_2 , 0 , buf_splitterfromN53_n129_1 );
buf_AQFP buf_splitterfromN56_n77_4_( clk_5 , splitterfromN56 , 0 , buf_splitterfromN56_n77_4 );
buf_AQFP buf_splitterfromN56_n77_3_( clk_7 , buf_splitterfromN56_n77_4 , 0 , buf_splitterfromN56_n77_3 );
buf_AQFP buf_splitterfromN56_n77_2_( clk_1 , buf_splitterfromN56_n77_3 , 0 , buf_splitterfromN56_n77_2 );
buf_AQFP buf_splitterfromN56_n77_1_( clk_3 , buf_splitterfromN56_n77_2 , 0 , buf_splitterfromN56_n77_1 );
buf_AQFP buf_splitterfromN60_n110_3_( clk_6 , splitterfromN60 , 0 , buf_splitterfromN60_n110_3 );
buf_AQFP buf_splitterfromN60_n110_2_( clk_8 , buf_splitterfromN60_n110_3 , 0 , buf_splitterfromN60_n110_2 );
buf_AQFP buf_splitterfromN60_n110_1_( clk_2 , buf_splitterfromN60_n110_2 , 0 , buf_splitterfromN60_n110_1 );
buf_AQFP buf_splitterfromN69_n79_3_( clk_4 , splitterfromN69 , 0 , buf_splitterfromN69_n79_3 );
buf_AQFP buf_splitterfromN69_n79_2_( clk_6 , buf_splitterfromN69_n79_3 , 0 , buf_splitterfromN69_n79_2 );
buf_AQFP buf_splitterfromN69_n79_1_( clk_8 , buf_splitterfromN69_n79_2 , 0 , buf_splitterfromN69_n79_1 );
buf_AQFP buf_splitterfromN73_n107_3_( clk_6 , splitterfromN73 , 0 , buf_splitterfromN73_n107_3 );
buf_AQFP buf_splitterfromN73_n107_2_( clk_8 , buf_splitterfromN73_n107_3 , 0 , buf_splitterfromN73_n107_2 );
buf_AQFP buf_splitterfromN73_n107_1_( clk_2 , buf_splitterfromN73_n107_2 , 0 , buf_splitterfromN73_n107_1 );
buf_AQFP buf_splitterfromN76_n57_3_( clk_5 , splitterfromN76 , 0 , buf_splitterfromN76_n57_3 );
buf_AQFP buf_splitterfromN76_n57_2_( clk_7 , buf_splitterfromN76_n57_3 , 0 , buf_splitterfromN76_n57_2 );
buf_AQFP buf_splitterfromN76_n57_1_( clk_1 , buf_splitterfromN76_n57_2 , 0 , buf_splitterfromN76_n57_1 );
buf_AQFP buf_splitterfromN79_n137_3_( clk_8 , splitterfromN79 , 0 , buf_splitterfromN79_n137_3 );
buf_AQFP buf_splitterfromN79_n137_2_( clk_2 , buf_splitterfromN79_n137_3 , 0 , buf_splitterfromN79_n137_2 );
buf_AQFP buf_splitterfromN79_n137_1_( clk_4 , buf_splitterfromN79_n137_2 , 0 , buf_splitterfromN79_n137_1 );
buf_AQFP buf_splitterfromN8_n100_3_( clk_7 , splitterfromN8 , 0 , buf_splitterfromN8_n100_3 );
buf_AQFP buf_splitterfromN8_n100_2_( clk_1 , buf_splitterfromN8_n100_3 , 0 , buf_splitterfromN8_n100_2 );
buf_AQFP buf_splitterfromN8_n100_1_( clk_3 , buf_splitterfromN8_n100_2 , 0 , buf_splitterfromN8_n100_1 );
buf_AQFP buf_splitterfromN82_n58_4_( clk_5 , splitterfromN82 , 0 , buf_splitterfromN82_n58_4 );
buf_AQFP buf_splitterfromN82_n58_3_( clk_7 , buf_splitterfromN82_n58_4 , 0 , buf_splitterfromN82_n58_3 );
buf_AQFP buf_splitterfromN82_n58_2_( clk_1 , buf_splitterfromN82_n58_3 , 0 , buf_splitterfromN82_n58_2 );
buf_AQFP buf_splitterfromN82_n58_1_( clk_3 , buf_splitterfromN82_n58_2 , 0 , buf_splitterfromN82_n58_1 );
buf_AQFP buf_splitterfromN86_n103_3_( clk_7 , splitterfromN86 , 0 , buf_splitterfromN86_n103_3 );
buf_AQFP buf_splitterfromN86_n103_2_( clk_1 , buf_splitterfromN86_n103_3 , 0 , buf_splitterfromN86_n103_2 );
buf_AQFP buf_splitterfromN86_n103_1_( clk_3 , buf_splitterfromN86_n103_2 , 0 , buf_splitterfromN86_n103_1 );
buf_AQFP buf_splitterfromN89_n72_3_( clk_5 , splitterfromN89 , 0 , buf_splitterfromN89_n72_3 );
buf_AQFP buf_splitterfromN89_n72_2_( clk_7 , buf_splitterfromN89_n72_3 , 0 , buf_splitterfromN89_n72_2 );
buf_AQFP buf_splitterfromN89_n72_1_( clk_1 , buf_splitterfromN89_n72_2 , 0 , buf_splitterfromN89_n72_1 );
buf_AQFP buf_splitterfromN92_n135_3_( clk_1 , splitterfromN92 , 0 , buf_splitterfromN92_n135_3 );
buf_AQFP buf_splitterfromN92_n135_2_( clk_3 , buf_splitterfromN92_n135_3 , 0 , buf_splitterfromN92_n135_2 );
buf_AQFP buf_splitterfromN92_n135_1_( clk_5 , buf_splitterfromN92_n135_2 , 0 , buf_splitterfromN92_n135_1 );
buf_AQFP buf_splitterfromN95_n73_4_( clk_5 , splitterfromN95 , 0 , buf_splitterfromN95_n73_4 );
buf_AQFP buf_splitterfromN95_n73_3_( clk_7 , buf_splitterfromN95_n73_4 , 0 , buf_splitterfromN95_n73_3 );
buf_AQFP buf_splitterfromN95_n73_2_( clk_1 , buf_splitterfromN95_n73_3 , 0 , buf_splitterfromN95_n73_2 );
buf_AQFP buf_splitterfromN95_n73_1_( clk_3 , buf_splitterfromN95_n73_2 , 0 , buf_splitterfromN95_n73_1 );
buf_AQFP buf_splitterfromN99_n92_2_( clk_7 , splitterfromN99 , 0 , buf_splitterfromN99_n92_2 );
buf_AQFP buf_splitterfromN99_n92_1_( clk_1 , buf_splitterfromN99_n92_2 , 0 , buf_splitterfromN99_n92_1 );
buf_AQFP buf_splitterfromn37_n62_2_( clk_8 , splitterfromn37 , 0 , buf_splitterfromn37_n62_2 );
buf_AQFP buf_splitterfromn37_n62_1_( clk_2 , buf_splitterfromn37_n62_2 , 0 , buf_splitterfromn37_n62_1 );
buf_AQFP buf_splitterfromn45_n80_3_( clk_6 , splitterfromn45 , 0 , buf_splitterfromn45_n80_3 );
buf_AQFP buf_splitterfromn45_n80_2_( clk_8 , buf_splitterfromn45_n80_3 , 0 , buf_splitterfromn45_n80_2 );
buf_AQFP buf_splitterfromn45_n80_1_( clk_2 , buf_splitterfromn45_n80_2 , 0 , buf_splitterfromn45_n80_1 );
buf_AQFP buf_splittern53ton69N223_N223_14_( clk_4 , splittern53ton69N223 , 0 , buf_splittern53ton69N223_N223_14 );
buf_AQFP buf_splittern53ton69N223_N223_13_( clk_6 , buf_splittern53ton69N223_N223_14 , 0 , buf_splittern53ton69N223_N223_13 );
buf_AQFP buf_splittern53ton69N223_N223_12_( clk_8 , buf_splittern53ton69N223_N223_13 , 0 , buf_splittern53ton69N223_N223_12 );
buf_AQFP buf_splittern53ton69N223_N223_11_( clk_2 , buf_splittern53ton69N223_N223_12 , 0 , buf_splittern53ton69N223_N223_11 );
buf_AQFP buf_splittern53ton69N223_N223_10_( clk_4 , buf_splittern53ton69N223_N223_11 , 0 , buf_splittern53ton69N223_N223_10 );
buf_AQFP buf_splittern53ton69N223_N223_9_( clk_6 , buf_splittern53ton69N223_N223_10 , 0 , buf_splittern53ton69N223_N223_9 );
buf_AQFP buf_splittern53ton69N223_N223_8_( clk_8 , buf_splittern53ton69N223_N223_9 , 0 , buf_splittern53ton69N223_N223_8 );
buf_AQFP buf_splittern53ton69N223_N223_7_( clk_2 , buf_splittern53ton69N223_N223_8 , 0 , buf_splittern53ton69N223_N223_7 );
buf_AQFP buf_splittern53ton69N223_N223_6_( clk_4 , buf_splittern53ton69N223_N223_7 , 0 , buf_splittern53ton69N223_N223_6 );
buf_AQFP buf_splittern53ton69N223_N223_5_( clk_6 , buf_splittern53ton69N223_N223_6 , 0 , buf_splittern53ton69N223_N223_5 );
buf_AQFP buf_splittern53ton69N223_N223_4_( clk_8 , buf_splittern53ton69N223_N223_5 , 0 , buf_splittern53ton69N223_N223_4 );
buf_AQFP buf_splittern53ton69N223_N223_3_( clk_2 , buf_splittern53ton69N223_N223_4 , 0 , buf_splittern53ton69N223_N223_3 );
buf_AQFP buf_splittern53ton69N223_N223_2_( clk_4 , buf_splittern53ton69N223_N223_3 , 0 , buf_splittern53ton69N223_N223_2 );
buf_AQFP buf_splittern53ton69N223_N223_1_( clk_6 , buf_splittern53ton69N223_N223_2 , 0 , buf_splittern53ton69N223_N223_1 );
buf_AQFP buf_splitterfromn55_n118_3_( clk_7 , splitterfromn55 , 0 , buf_splitterfromn55_n118_3 );
buf_AQFP buf_splitterfromn55_n118_2_( clk_1 , buf_splitterfromn55_n118_3 , 0 , buf_splitterfromn55_n118_2 );
buf_AQFP buf_splitterfromn55_n118_1_( clk_3 , buf_splitterfromn55_n118_2 , 0 , buf_splitterfromn55_n118_1 );
buf_AQFP buf_splitterfromn58_n104_3_( clk_7 , splitterfromn58 , 0 , buf_splitterfromn58_n104_3 );
buf_AQFP buf_splitterfromn58_n104_2_( clk_1 , buf_splitterfromn58_n104_3 , 0 , buf_splitterfromn58_n104_2 );
buf_AQFP buf_splitterfromn58_n104_1_( clk_3 , buf_splitterfromn58_n104_2 , 0 , buf_splitterfromn58_n104_1 );
buf_AQFP buf_splitterfromn62_n90_3_( clk_7 , splitterfromn62 , 0 , buf_splitterfromn62_n90_3 );
buf_AQFP buf_splitterfromn62_n90_2_( clk_1 , buf_splitterfromn62_n90_3 , 0 , buf_splitterfromn62_n90_2 );
buf_AQFP buf_splitterfromn62_n90_1_( clk_3 , buf_splitterfromn62_n90_2 , 0 , buf_splitterfromn62_n90_1 );
buf_AQFP buf_splitterfromn65_n96_3_( clk_7 , splitterfromn65 , 0 , buf_splitterfromn65_n96_3 );
buf_AQFP buf_splitterfromn65_n96_2_( clk_1 , buf_splitterfromn65_n96_3 , 0 , buf_splitterfromn65_n96_2 );
buf_AQFP buf_splitterfromn65_n96_1_( clk_3 , buf_splitterfromn65_n96_2 , 0 , buf_splitterfromn65_n96_1 );
buf_AQFP buf_splitterfromn70_n101_3_( clk_7 , splitterfromn70 , 0 , buf_splitterfromn70_n101_3 );
buf_AQFP buf_splitterfromn70_n101_2_( clk_1 , buf_splitterfromn70_n101_3 , 0 , buf_splitterfromn70_n101_2 );
buf_AQFP buf_splitterfromn70_n101_1_( clk_3 , buf_splitterfromn70_n101_2 , 0 , buf_splitterfromn70_n101_1 );
buf_AQFP buf_splitterfromn73_n93_3_( clk_7 , splitterfromn73 , 0 , buf_splitterfromn73_n93_3 );
buf_AQFP buf_splitterfromn73_n93_2_( clk_1 , buf_splitterfromn73_n93_3 , 0 , buf_splitterfromn73_n93_2 );
buf_AQFP buf_splitterfromn73_n93_1_( clk_3 , buf_splitterfromn73_n93_2 , 0 , buf_splitterfromn73_n93_1 );
buf_AQFP buf_splitterfromn77_n111_3_( clk_7 , splitterfromn77 , 0 , buf_splitterfromn77_n111_3 );
buf_AQFP buf_splitterfromn77_n111_2_( clk_1 , buf_splitterfromn77_n111_3 , 0 , buf_splitterfromn77_n111_2 );
buf_AQFP buf_splitterfromn77_n111_1_( clk_3 , buf_splitterfromn77_n111_2 , 0 , buf_splitterfromn77_n111_1 );
buf_AQFP buf_splitterfromn80_n108_4_( clk_6 , splitterfromn80 , 0 , buf_splitterfromn80_n108_4 );
buf_AQFP buf_splitterfromn80_n108_3_( clk_8 , buf_splitterfromn80_n108_4 , 0 , buf_splitterfromn80_n108_3 );
buf_AQFP buf_splitterfromn80_n108_2_( clk_2 , buf_splitterfromn80_n108_3 , 0 , buf_splitterfromn80_n108_2 );
buf_AQFP buf_splitterfromn80_n108_1_( clk_4 , buf_splitterfromn80_n108_2 , 0 , buf_splitterfromn80_n108_1 );
buf_AQFP buf_splitterfromn83_n115_4_( clk_6 , splitterfromn83 , 0 , buf_splitterfromn83_n115_4 );
buf_AQFP buf_splitterfromn83_n115_3_( clk_8 , buf_splitterfromn83_n115_4 , 0 , buf_splitterfromn83_n115_3 );
buf_AQFP buf_splitterfromn83_n115_2_( clk_2 , buf_splitterfromn83_n115_3 , 0 , buf_splitterfromn83_n115_2 );
buf_AQFP buf_splitterfromn83_n115_1_( clk_4 , buf_splitterfromn83_n115_2 , 0 , buf_splitterfromn83_n115_1 );
buf_AQFP buf_splittern88ton117N329_N329_9_( clk_5 , splittern88ton117N329 , 0 , buf_splittern88ton117N329_N329_9 );
buf_AQFP buf_splittern88ton117N329_N329_8_( clk_7 , buf_splittern88ton117N329_N329_9 , 0 , buf_splittern88ton117N329_N329_8 );
buf_AQFP buf_splittern88ton117N329_N329_7_( clk_1 , buf_splittern88ton117N329_N329_8 , 0 , buf_splittern88ton117N329_N329_7 );
buf_AQFP buf_splittern88ton117N329_N329_6_( clk_3 , buf_splittern88ton117N329_N329_7 , 0 , buf_splittern88ton117N329_N329_6 );
buf_AQFP buf_splittern88ton117N329_N329_5_( clk_5 , buf_splittern88ton117N329_N329_6 , 0 , buf_splittern88ton117N329_N329_5 );
buf_AQFP buf_splittern88ton117N329_N329_4_( clk_7 , buf_splittern88ton117N329_N329_5 , 0 , buf_splittern88ton117N329_N329_4 );
buf_AQFP buf_splittern88ton117N329_N329_3_( clk_1 , buf_splittern88ton117N329_N329_4 , 0 , buf_splittern88ton117N329_N329_3 );
buf_AQFP buf_splittern88ton117N329_N329_2_( clk_3 , buf_splittern88ton117N329_N329_3 , 0 , buf_splittern88ton117N329_N329_2 );
buf_AQFP buf_splittern88ton117N329_N329_1_( clk_5 , buf_splittern88ton117N329_N329_2 , 0 , buf_splittern88ton117N329_N329_1 );
buf_AQFP buf_splitterfromn90_n125_3_( clk_1 , splitterfromn90 , 0 , buf_splitterfromn90_n125_3 );
buf_AQFP buf_splitterfromn90_n125_2_( clk_3 , buf_splitterfromn90_n125_3 , 0 , buf_splitterfromn90_n125_2 );
buf_AQFP buf_splitterfromn90_n125_1_( clk_5 , buf_splitterfromn90_n125_2 , 0 , buf_splitterfromn90_n125_1 );
buf_AQFP buf_splitterfromn93_n141_3_( clk_1 , splitterfromn93 , 0 , buf_splitterfromn93_n141_3 );
buf_AQFP buf_splitterfromn93_n141_2_( clk_3 , buf_splitterfromn93_n141_3 , 0 , buf_splitterfromn93_n141_2 );
buf_AQFP buf_splitterfromn93_n141_1_( clk_5 , buf_splitterfromn93_n141_2 , 0 , buf_splitterfromn93_n141_1 );
buf_AQFP buf_splitterfromn96_n127_3_( clk_1 , splitterfromn96 , 0 , buf_splitterfromn96_n127_3 );
buf_AQFP buf_splitterfromn96_n127_2_( clk_3 , buf_splitterfromn96_n127_3 , 0 , buf_splitterfromn96_n127_2 );
buf_AQFP buf_splitterfromn96_n127_1_( clk_5 , buf_splitterfromn96_n127_2 , 0 , buf_splitterfromn96_n127_1 );
buf_AQFP buf_splitterfromn101_n148_4_( clk_1 , splitterfromn101 , 0 , buf_splitterfromn101_n148_4 );
buf_AQFP buf_splitterfromn101_n148_3_( clk_3 , buf_splitterfromn101_n148_4 , 0 , buf_splitterfromn101_n148_3 );
buf_AQFP buf_splitterfromn101_n148_2_( clk_5 , buf_splitterfromn101_n148_3 , 0 , buf_splitterfromn101_n148_2 );
buf_AQFP buf_splitterfromn101_n148_1_( clk_7 , buf_splitterfromn101_n148_2 , 0 , buf_splitterfromn101_n148_1 );
buf_AQFP buf_splitterfromn104_n136_3_( clk_1 , splitterfromn104 , 0 , buf_splitterfromn104_n136_3 );
buf_AQFP buf_splitterfromn104_n136_2_( clk_3 , buf_splitterfromn104_n136_3 , 0 , buf_splitterfromn104_n136_2 );
buf_AQFP buf_splitterfromn104_n136_1_( clk_5 , buf_splitterfromn104_n136_2 , 0 , buf_splitterfromn104_n136_1 );
buf_AQFP buf_splitterfromn108_n138_4_( clk_8 , splitterfromn108 , 0 , buf_splitterfromn108_n138_4 );
buf_AQFP buf_splitterfromn108_n138_3_( clk_2 , buf_splitterfromn108_n138_4 , 0 , buf_splitterfromn108_n138_3 );
buf_AQFP buf_splitterfromn108_n138_2_( clk_4 , buf_splitterfromn108_n138_3 , 0 , buf_splitterfromn108_n138_2 );
buf_AQFP buf_splitterfromn108_n138_1_( clk_6 , buf_splitterfromn108_n138_2 , 0 , buf_splitterfromn108_n138_1 );
buf_AQFP buf_splitterfromn111_n131_4_( clk_7 , splitterfromn111 , 0 , buf_splitterfromn111_n131_4 );
buf_AQFP buf_splitterfromn111_n131_3_( clk_1 , buf_splitterfromn111_n131_4 , 0 , buf_splitterfromn111_n131_3 );
buf_AQFP buf_splitterfromn111_n131_2_( clk_3 , buf_splitterfromn111_n131_3 , 0 , buf_splitterfromn111_n131_2 );
buf_AQFP buf_splitterfromn111_n131_1_( clk_5 , buf_splitterfromn111_n131_2 , 0 , buf_splitterfromn111_n131_1 );
buf_AQFP buf_splitterfromn112_n132_3_( clk_1 , splitterfromn112 , 0 , buf_splitterfromn112_n132_3 );
buf_AQFP buf_splitterfromn112_n132_2_( clk_3 , buf_splitterfromn112_n132_3 , 0 , buf_splitterfromn112_n132_2 );
buf_AQFP buf_splitterfromn112_n132_1_( clk_5 , buf_splitterfromn112_n132_2 , 0 , buf_splitterfromn112_n132_1 );
buf_AQFP buf_splitterfromn115_n130_4_( clk_8 , splitterfromn115 , 0 , buf_splitterfromn115_n130_4 );
buf_AQFP buf_splitterfromn115_n130_3_( clk_2 , buf_splitterfromn115_n130_4 , 0 , buf_splitterfromn115_n130_3 );
buf_AQFP buf_splitterfromn115_n130_2_( clk_4 , buf_splitterfromn115_n130_3 , 0 , buf_splitterfromn115_n130_2 );
buf_AQFP buf_splitterfromn115_n130_1_( clk_6 , buf_splitterfromn115_n130_2 , 0 , buf_splitterfromn115_n130_1 );
buf_AQFP buf_splitterfromn118_n143_4_( clk_8 , splitterfromn118 , 0 , buf_splitterfromn118_n143_4 );
buf_AQFP buf_splitterfromn118_n143_3_( clk_2 , buf_splitterfromn118_n143_4 , 0 , buf_splitterfromn118_n143_3 );
buf_AQFP buf_splitterfromn118_n143_2_( clk_4 , buf_splitterfromn118_n143_3 , 0 , buf_splitterfromn118_n143_2 );
buf_AQFP buf_splitterfromn118_n143_1_( clk_6 , buf_splitterfromn118_n143_2 , 0 , buf_splitterfromn118_n143_1 );
buf_AQFP buf_splittern123ton140N370_N370_4_( clk_7 , splittern123ton140N370 , 0 , buf_splittern123ton140N370_N370_4 );
buf_AQFP buf_splittern123ton140N370_N370_3_( clk_1 , buf_splittern123ton140N370_N370_4 , 0 , buf_splittern123ton140N370_N370_3 );
buf_AQFP buf_splittern123ton140N370_N370_2_( clk_3 , buf_splittern123ton140N370_N370_3 , 0 , buf_splittern123ton140N370_N370_2 );
buf_AQFP buf_splittern123ton140N370_N370_1_( clk_5 , buf_splittern123ton140N370_N370_2 , 0 , buf_splittern123ton140N370_N370_1 );
buf_AQFP buf_splitterfromn125_n156_2_( clk_2 , splitterfromn125 , 0 , buf_splitterfromn125_n156_2 );
buf_AQFP buf_splitterfromn125_n156_1_( clk_4 , buf_splitterfromn125_n156_2 , 0 , buf_splitterfromn125_n156_1 );
buf_AQFP buf_splitterfromn127_n157_2_( clk_2 , splitterfromn127 , 0 , buf_splitterfromn127_n157_2 );
buf_AQFP buf_splitterfromn127_n157_1_( clk_4 , buf_splitterfromn127_n157_2 , 0 , buf_splitterfromn127_n157_1 );
buf_AQFP buf_splitterfromn134_N430_1_( clk_6 , splitterfromn134 , 0 , buf_splitterfromn134_N430_1 );
buf_AQFP buf_splitterfromn138_n152_1_( clk_2 , splitterfromn138 , 0 , buf_splitterfromn138_n152_1 );
splitter_AQFP splitterfromN1_( clk_3 , N1 , 0 , splitterfromN1 );
splitter_AQFP splitterfromN102_( clk_5 , buf_N102_splitterfromN102_1 , 0 , splitterfromN102 );
splitter_AQFP splitterfromN105_( clk_7 , buf_N105_splitterfromN105_1 , 0 , splitterfromN105 );
splitter_AQFP splitterfromN108_( clk_5 , buf_N108_splitterfromN108_1 , 0 , splitterfromN108 );
splitter_AQFP splitterfromN11_( clk_3 , N11 , 0 , splitterfromN11 );
splitter_AQFP splitterfromN112_( clk_4 , buf_N112_splitterfromN112_1 , 0 , splitterfromN112 );
splitter_AQFP splitterfromN115_( clk_6 , buf_N115_splitterfromN115_1 , 0 , splitterfromN115 );
splitter_AQFP splitterfromN14_( clk_7 , buf_N14_splitterfromN14_1 , 0 , splitterfromN14 );
splitter_AQFP splitterfromN17_( clk_3 , N17 , 0 , splitterfromN17 );
splitter_AQFP splitterfromN21_( clk_5 , buf_N21_splitterfromN21_1 , 0 , splitterfromN21 );
splitter_AQFP splitterfromN27_( clk_7 , buf_N27_splitterfromN27_1 , 0 , splitterfromN27 );
splitter_AQFP splitterfromN30_( clk_3 , N30 , 0 , splitterfromN30 );
splitter_AQFP splitterfromN34_( clk_5 , buf_N34_splitterfromN34_1 , 0 , splitterfromN34 );
splitter_AQFP splitterfromN37_( clk_3 , N37 , 0 , splitterfromN37 );
splitter_AQFP splitterfromN4_( clk_4 , buf_N4_splitterfromN4_1 , 0 , splitterfromN4 );
splitter_AQFP splitterfromN40_( clk_7 , buf_N40_splitterfromN40_1 , 0 , splitterfromN40 );
splitter_AQFP splitterfromN43_( clk_3 , N43 , 0 , splitterfromN43 );
splitter_AQFP splitterfromN47_( clk_4 , buf_N47_splitterfromN47_1 , 0 , splitterfromN47 );
splitter_AQFP splitterfromN50_( clk_3 , N50 , 0 , splitterfromN50 );
splitter_AQFP splitterfromN53_( clk_6 , buf_N53_splitterfromN53_1 , 0 , splitterfromN53 );
splitter_AQFP splitterfromN56_( clk_3 , N56 , 0 , splitterfromN56 );
splitter_AQFP splitterfromN60_( clk_4 , buf_N60_splitterfromN60_1 , 0 , splitterfromN60 );
splitter_AQFP splitterfromN69_( clk_2 , N69 , 0 , splitterfromN69 );
splitter_AQFP splitterfromN73_( clk_4 , buf_N73_splitterfromN73_1 , 0 , splitterfromN73 );
splitter_AQFP splitterfromN76_( clk_3 , N76 , 0 , splitterfromN76 );
splitter_AQFP splitterfromN79_( clk_6 , buf_N79_splitterfromN79_1 , 0 , splitterfromN79 );
splitter_AQFP splitterfromN8_( clk_5 , buf_N8_splitterfromN8_1 , 0 , splitterfromN8 );
splitter_AQFP splitterfromN82_( clk_3 , N82 , 0 , splitterfromN82 );
splitter_AQFP splitterfromN86_( clk_5 , buf_N86_splitterfromN86_1 , 0 , splitterfromN86 );
splitter_AQFP splitterfromN89_( clk_3 , N89 , 0 , splitterfromN89 );
splitter_AQFP splitterfromN92_( clk_7 , buf_N92_splitterfromN92_1 , 0 , splitterfromN92 );
splitter_AQFP splitterfromN95_( clk_3 , N95 , 0 , splitterfromN95 );
splitter_AQFP splitterfromN99_( clk_5 , buf_N99_splitterfromN99_1 , 0 , splitterfromN99 );
splitter_AQFP splitterfromn37_( clk_6 , n37 , 0 , splitterfromn37 );
splitter_AQFP splitterfromn45_( clk_4 , n45 , 0 , splitterfromn45 );
splitter_AQFP splittern53ton79N223_( clk_1 , n53 , 0 , splittern53ton79N223 );
splitter_AQFP splittern53ton54n64_( clk_2 , splittern53ton79N223 , 0 , splittern53ton54n64 );
splitter_AQFP splittern53ton69N223_( clk_2 , splittern53ton79N223 , 0 , splittern53ton69N223 );
splitter_AQFP splitterfromn55_( clk_5 , n55 , 0 , splitterfromn55 );
splitter_AQFP splitterfromn58_( clk_5 , n58 , 0 , splitterfromn58 );
splitter_AQFP splitterfromn62_( clk_5 , n62 , 0 , splitterfromn62 );
splitter_AQFP splitterfromn65_( clk_5 , n65 , 0 , splitterfromn65 );
splitter_AQFP splitterfromn70_( clk_5 , n70 , 0 , splitterfromn70 );
splitter_AQFP splitterfromn73_( clk_5 , n73 , 0 , splitterfromn73 );
splitter_AQFP splitterfromn77_( clk_5 , n77 , 0 , splitterfromn77 );
splitter_AQFP splitterfromn80_( clk_4 , n80 , 0 , splitterfromn80 );
splitter_AQFP splitterfromn83_( clk_4 , n83 , 0 , splitterfromn83 );
splitter_AQFP splittern88ton110N329_( clk_2 , n88 , 0 , splittern88ton110N329 );
splitter_AQFP splittern88ton100n114_( clk_3 , splittern88ton110N329 , 0 , splittern88ton100n114 );
splitter_AQFP splittern88ton117N329_( clk_3 , splittern88ton110N329 , 0 , splittern88ton117N329 );
splitter_AQFP splitterfromn90_( clk_7 , n90 , 0 , splitterfromn90 );
splitter_AQFP splitterfromn93_( clk_7 , n93 , 0 , splitterfromn93 );
splitter_AQFP splitterfromn96_( clk_7 , n96 , 0 , splitterfromn96 );
splitter_AQFP splitterfromn101_( clk_7 , n101 , 0 , splitterfromn101 );
splitter_AQFP splitterfromn104_( clk_7 , n104 , 0 , splitterfromn104 );
splitter_AQFP splitterfromn108_( clk_6 , n108 , 0 , splitterfromn108 );
splitter_AQFP splitterfromn111_( clk_5 , n111 , 0 , splitterfromn111 );
splitter_AQFP splitterfromn112_( clk_7 , n112 , 0 , splitterfromn112 );
splitter_AQFP splitterfromn115_( clk_6 , n115 , 0 , splitterfromn115 );
splitter_AQFP splitterfromn118_( clk_6 , n118 , 0 , splitterfromn118 );
splitter_AQFP splittern123ton124N370_( clk_4 , n123 , 0 , splittern123ton124N370 );
splitter_AQFP splittern123ton129n137_( clk_5 , splittern123ton124N370 , 0 , splittern123ton129n137 );
splitter_AQFP splittern123ton140N370_( clk_5 , splittern123ton124N370 , 0 , splittern123ton140N370 );
splitter_AQFP splitterfromn125_( clk_8 , n125 , 0 , splitterfromn125 );
splitter_AQFP splitterfromn127_( clk_8 , n127 , 0 , splitterfromn127 );
splitter_AQFP splitterfromn128_( clk_2 , n128 , 0 , splitterfromn128 );
splitter_AQFP splitterfromn130_( clk_8 , n130 , 0 , splitterfromn130 );
splitter_AQFP splittern133ton134n152_( clk_2 , n133 , 0 , splittern133ton134n152 );
splitter_AQFP splitterfromn134_( clk_4 , n134 , 0 , splitterfromn134 );
splitter_AQFP splitterfromn136_( clk_8 , n136 , 0 , splitterfromn136 );
splitter_AQFP splitterfromn138_( clk_8 , n138 , 0 , splitterfromn138 );
splitter_AQFP splitterfromn139_( clk_2 , n139 , 0 , splitterfromn139 );
splitter_AQFP splitterfromn141_( clk_8 , n141 , 0 , splitterfromn141 );

endmodule