module top( clk_1 , clk_2 , clk_3 , clk_4 , clk_5 , clk_6 , clk_7 , clk_8 , G1 , G10 , G100 , G101 , G102 , G103 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 , G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2591 , G2593 , G2594 );

input G1 , G10 , G100 , G101 , G102 , G103 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 ;
output G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2591 , G2593 , G2594 ;
wire n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , buf_G10_splitterfromG10_11 , buf_G10_splitterfromG10_10 , buf_G10_splitterfromG10_9 , buf_G10_splitterfromG10_8 , buf_G10_splitterfromG10_7 , buf_G10_splitterfromG10_6 , buf_G10_splitterfromG10_5 , buf_G10_splitterfromG10_4 , buf_G10_splitterfromG10_3 , buf_G10_splitterfromG10_2 , buf_G10_splitterfromG10_1 , buf_G100_n195_1 , buf_G101_n388_2 , buf_G101_n388_1 , buf_G102_n373_2 , buf_G102_n373_1 , buf_G103_n354_2 , buf_G103_n354_1 , buf_G105_n304_2 , buf_G105_n304_1 , buf_G106_splitterfromG106_7 , buf_G106_splitterfromG106_6 , buf_G106_splitterfromG106_5 , buf_G106_splitterfromG106_4 , buf_G106_splitterfromG106_3 , buf_G106_splitterfromG106_2 , buf_G106_splitterfromG106_1 , buf_G107_n291_2 , buf_G107_n291_1 , buf_G108_n185_2 , buf_G108_n185_1 , buf_G109_n178_1 , buf_G11_n162_1 , buf_G110_n196_1 , buf_G111_n390_2 , buf_G111_n390_1 , buf_G112_n375_2 , buf_G112_n375_1 , buf_G113_n356_2 , buf_G113_n356_1 , buf_G116_n233_1 , buf_G118_splitterfromG118_5 , buf_G118_splitterfromG118_4 , buf_G118_splitterfromG118_3 , buf_G118_splitterfromG118_2 , buf_G118_splitterfromG118_1 , buf_G119_splitterfromG119_9 , buf_G119_splitterfromG119_8 , buf_G119_splitterfromG119_7 , buf_G119_splitterfromG119_6 , buf_G119_splitterfromG119_5 , buf_G119_splitterfromG119_4 , buf_G119_splitterfromG119_3 , buf_G119_splitterfromG119_2 , buf_G119_splitterfromG119_1 , buf_G122_splitterG122ton437n438_6 , buf_G122_splitterG122ton437n438_5 , buf_G122_splitterG122ton437n438_4 , buf_G122_splitterG122ton437n438_3 , buf_G122_splitterG122ton437n438_2 , buf_G122_splitterG122ton437n438_1 , buf_G123_splitterG123ton285n447_5 , buf_G123_splitterG123ton285n447_4 , buf_G123_splitterG123ton285n447_3 , buf_G123_splitterG123ton285n447_2 , buf_G123_splitterG123ton285n447_1 , buf_G124_splitterfromG124_13 , buf_G124_splitterfromG124_12 , buf_G124_splitterfromG124_11 , buf_G124_splitterfromG124_10 , buf_G124_splitterfromG124_9 , buf_G124_splitterfromG124_8 , buf_G124_splitterfromG124_7 , buf_G124_splitterfromG124_6 , buf_G124_splitterfromG124_5 , buf_G124_splitterfromG124_4 , buf_G124_splitterfromG124_3 , buf_G124_splitterfromG124_2 , buf_G124_splitterfromG124_1 , buf_G125_splitterfromG125_5 , buf_G125_splitterfromG125_4 , buf_G125_splitterfromG125_3 , buf_G125_splitterfromG125_2 , buf_G125_splitterfromG125_1 , buf_G126_splitterfromG126_4 , buf_G126_splitterfromG126_3 , buf_G126_splitterfromG126_2 , buf_G126_splitterfromG126_1 , buf_G127_n448_3 , buf_G127_n448_2 , buf_G127_n448_1 , buf_G128_splitterfromG128_4 , buf_G128_splitterfromG128_3 , buf_G128_splitterfromG128_2 , buf_G128_splitterfromG128_1 , buf_G129_splitterfromG129_4 , buf_G129_splitterfromG129_3 , buf_G129_splitterfromG129_2 , buf_G129_splitterfromG129_1 , buf_G130_splitterfromG130_4 , buf_G130_splitterfromG130_3 , buf_G130_splitterfromG130_2 , buf_G130_splitterfromG130_1 , buf_G131_splitterG131ton368n487_5 , buf_G131_splitterG131ton368n487_4 , buf_G131_splitterG131ton368n487_3 , buf_G131_splitterG131ton368n487_2 , buf_G131_splitterG131ton368n487_1 , buf_G132_splitterfromG132_5 , buf_G132_splitterfromG132_4 , buf_G132_splitterfromG132_3 , buf_G132_splitterfromG132_2 , buf_G132_splitterfromG132_1 , buf_G133_splitterfromG133_5 , buf_G133_splitterfromG133_4 , buf_G133_splitterfromG133_3 , buf_G133_splitterfromG133_2 , buf_G133_splitterfromG133_1 , buf_G134_splitterG134ton513n401_3 , buf_G134_splitterG134ton513n401_2 , buf_G134_splitterG134ton513n401_1 , buf_G135_splitterG135ton505n309_3 , buf_G135_splitterG135ton505n309_2 , buf_G135_splitterG135ton505n309_1 , buf_G136_splitterG136ton500n469_3 , buf_G136_splitterG136ton500n469_2 , buf_G136_splitterG136ton500n469_1 , buf_G137_splitterG137toG2536G2538_13 , buf_G137_splitterG137toG2536G2538_12 , buf_G137_splitterG137toG2536G2538_11 , buf_G137_splitterG137toG2536G2538_10 , buf_G137_splitterG137toG2536G2538_9 , buf_G137_splitterG137toG2536G2538_8 , buf_G137_splitterG137toG2536G2538_7 , buf_G137_splitterG137toG2536G2538_6 , buf_G137_splitterG137toG2536G2538_5 , buf_G137_splitterG137toG2536G2538_4 , buf_G137_splitterG137toG2536G2538_3 , buf_G137_splitterG137toG2536G2538_2 , buf_G137_splitterG137toG2536G2538_1 , buf_G138_splitterG138ton502n465_4 , buf_G138_splitterG138ton502n465_3 , buf_G138_splitterG138ton502n465_2 , buf_G138_splitterG138ton502n465_1 , buf_G139_splitterG139ton159n461_3 , buf_G139_splitterG139ton159n461_2 , buf_G139_splitterG139ton159n461_1 , buf_G14_n335_2 , buf_G14_n335_1 , buf_G140_splitterG140ton159n457_3 , buf_G140_splitterG140ton159n457_2 , buf_G140_splitterG140ton159n457_1 , buf_G141_splitterG141ton158n481_4 , buf_G141_splitterG141ton158n481_3 , buf_G141_splitterG141ton158n481_2 , buf_G141_splitterG141ton158n481_1 , buf_G142_splitterG142ton158n488_3 , buf_G142_splitterG142ton158n488_2 , buf_G142_splitterG142ton158n488_1 , buf_G143_splitterfromG143_3 , buf_G143_splitterfromG143_2 , buf_G143_splitterfromG143_1 , buf_G144_n298_5 , buf_G144_n298_4 , buf_G144_n298_3 , buf_G144_n298_2 , buf_G144_n298_1 , buf_G147_splitterfromG147_9 , buf_G147_splitterfromG147_8 , buf_G147_splitterfromG147_7 , buf_G147_splitterfromG147_6 , buf_G147_splitterfromG147_5 , buf_G147_splitterfromG147_4 , buf_G147_splitterfromG147_3 , buf_G147_splitterfromG147_2 , buf_G147_splitterfromG147_1 , buf_G15_n314_1 , buf_G16_n365_3 , buf_G16_n365_2 , buf_G16_n365_1 , buf_G17_n420_2 , buf_G17_n420_1 , buf_G18_n398_2 , buf_G18_n398_1 , buf_G19_n299_2 , buf_G19_n299_1 , buf_G20_n371_4 , buf_G20_n371_3 , buf_G20_n371_2 , buf_G20_n371_1 , buf_G21_n324_2 , buf_G21_n324_1 , buf_G24_n352_1 , buf_G25_n386_1 , buf_G26_n344_3 , buf_G26_n344_2 , buf_G26_n344_1 , buf_G27_n329_2 , buf_G27_n329_1 , buf_G28_n235_13 , buf_G28_n235_12 , buf_G28_n235_11 , buf_G28_n235_10 , buf_G28_n235_9 , buf_G28_n235_8 , buf_G28_n235_7 , buf_G28_n235_6 , buf_G28_n235_5 , buf_G28_n235_4 , buf_G28_n235_3 , buf_G28_n235_2 , buf_G28_n235_1 , buf_G29_n445_7 , buf_G29_n445_6 , buf_G29_n445_5 , buf_G29_n445_4 , buf_G29_n445_3 , buf_G29_n445_2 , buf_G29_n445_1 , buf_G30_n449_3 , buf_G30_n449_2 , buf_G30_n449_1 , buf_G31_n224_2 , buf_G31_n224_1 , buf_G32_splitterfromG32_7 , buf_G32_splitterfromG32_6 , buf_G32_splitterfromG32_5 , buf_G32_splitterfromG32_4 , buf_G32_splitterfromG32_3 , buf_G32_splitterfromG32_2 , buf_G32_splitterfromG32_1 , buf_G33_n260_1 , buf_G34_n252_1 , buf_G35_n247_2 , buf_G35_n247_1 , buf_G36_n199_1 , buf_G37_n208_1 , buf_G38_n216_1 , buf_G39_n238_1 , buf_G40_n268_1 , buf_G41_n429_2 , buf_G41_n429_1 , buf_G42_n228_2 , buf_G42_n228_1 , buf_G43_splitterfromG43_6 , buf_G43_splitterfromG43_5 , buf_G43_splitterfromG43_4 , buf_G43_splitterfromG43_3 , buf_G43_splitterfromG43_2 , buf_G43_splitterfromG43_1 , buf_G44_n264_2 , buf_G44_n264_1 , buf_G45_n256_2 , buf_G45_n256_1 , buf_G46_n204_1 , buf_G47_n212_2 , buf_G47_n212_1 , buf_G48_n220_2 , buf_G48_n220_1 , buf_G49_n242_2 , buf_G49_n242_1 , buf_G5_n320_1 , buf_G50_n272_2 , buf_G50_n272_1 , buf_G51_n433_2 , buf_G51_n433_1 , buf_G52_n229_2 , buf_G52_n229_1 , buf_G53_splitterfromG53_6 , buf_G53_splitterfromG53_5 , buf_G53_splitterfromG53_4 , buf_G53_splitterfromG53_3 , buf_G53_splitterfromG53_2 , buf_G53_splitterfromG53_1 , buf_G54_n265_2 , buf_G54_n265_1 , buf_G55_n257_2 , buf_G55_n257_1 , buf_G56_n246_2 , buf_G56_n246_1 , buf_G57_n205_2 , buf_G57_n205_1 , buf_G58_n213_2 , buf_G58_n213_1 , buf_G59_n221_2 , buf_G59_n221_1 , buf_G6_n404_3 , buf_G6_n404_2 , buf_G6_n404_1 , buf_G60_n243_2 , buf_G60_n243_1 , buf_G61_n273_2 , buf_G61_n273_1 , buf_G62_n434_2 , buf_G62_n434_1 , buf_G63_n225_1 , buf_G64_splitterfromG64_6 , buf_G64_splitterfromG64_5 , buf_G64_splitterfromG64_4 , buf_G64_splitterfromG64_3 , buf_G64_splitterfromG64_2 , buf_G64_splitterfromG64_1 , buf_G66_n253_1 , buf_G67_n248_1 , buf_G68_n200_1 , buf_G69_n209_1 , buf_G70_n217_1 , buf_G71_n239_1 , buf_G72_n269_1 , buf_G73_n430_1 , buf_G74_n163_1 , buf_G75_n300_2 , buf_G75_n300_1 , buf_G76_splitterfromG76_6 , buf_G76_splitterfromG76_5 , buf_G76_splitterfromG76_4 , buf_G76_splitterfromG76_3 , buf_G76_splitterfromG76_2 , buf_G76_splitterfromG76_1 , buf_G77_n288_2 , buf_G77_n288_1 , buf_G78_n189_2 , buf_G78_n189_1 , buf_G79_n179_1 , buf_G8_splitterG8ton451n486_5 , buf_G8_splitterG8ton451n486_4 , buf_G8_splitterG8ton451n486_3 , buf_G8_splitterG8ton451n486_2 , buf_G8_splitterG8ton451n486_1 , buf_G80_n192_1 , buf_G81_n387_2 , buf_G81_n387_1 , buf_G82_n372_2 , buf_G82_n372_1 , buf_G83_n357_2 , buf_G83_n357_1 , buf_G85_n301_2 , buf_G85_n301_1 , buf_G86_splitterfromG86_7 , buf_G86_splitterfromG86_6 , buf_G86_splitterfromG86_5 , buf_G86_splitterfromG86_4 , buf_G86_splitterfromG86_3 , buf_G86_splitterfromG86_2 , buf_G86_splitterfromG86_1 , buf_G87_n292_2 , buf_G87_n292_1 , buf_G88_n188_2 , buf_G88_n188_1 , buf_G89_n181_1 , buf_G9_n410_1 , buf_G90_n193_1 , buf_G91_n391_2 , buf_G91_n391_1 , buf_G92_n376_2 , buf_G92_n376_1 , buf_G93_n353_2 , buf_G93_n353_1 , buf_G95_n303_2 , buf_G95_n303_1 , buf_G96_splitterfromG96_7 , buf_G96_splitterfromG96_6 , buf_G96_splitterfromG96_5 , buf_G96_splitterfromG96_4 , buf_G96_splitterfromG96_3 , buf_G96_splitterfromG96_2 , buf_G96_splitterfromG96_1 , buf_G97_n289_2 , buf_G97_n289_1 , buf_G98_n186_2 , buf_G98_n186_1 , buf_G99_n182_1 , buf_n160_G2547_8 , buf_n160_G2547_7 , buf_n160_G2547_6 , buf_n160_G2547_5 , buf_n160_G2547_4 , buf_n160_G2547_3 , buf_n160_G2547_2 , buf_n160_G2547_1 , buf_n162_G2548_12 , buf_n162_G2548_11 , buf_n162_G2548_10 , buf_n162_G2548_9 , buf_n162_G2548_8 , buf_n162_G2548_7 , buf_n162_G2548_6 , buf_n162_G2548_5 , buf_n162_G2548_4 , buf_n162_G2548_3 , buf_n162_G2548_2 , buf_n162_G2548_1 , buf_n163_G2550_12 , buf_n163_G2550_11 , buf_n163_G2550_10 , buf_n163_G2550_9 , buf_n163_G2550_8 , buf_n163_G2550_7 , buf_n163_G2550_6 , buf_n163_G2550_5 , buf_n163_G2550_4 , buf_n163_G2550_3 , buf_n163_G2550_2 , buf_n163_G2550_1 , buf_n164_splittern164ton165G2551_8 , buf_n164_splittern164ton165G2551_7 , buf_n164_splittern164ton165G2551_6 , buf_n164_splittern164ton165G2551_5 , buf_n164_splittern164ton165G2551_4 , buf_n164_splittern164ton165G2551_3 , buf_n164_splittern164ton165G2551_2 , buf_n164_splittern164ton165G2551_1 , buf_n165_G2552_3 , buf_n165_G2552_2 , buf_n165_G2552_1 , buf_n166_G2553_3 , buf_n166_G2553_2 , buf_n166_G2553_1 , buf_n173_splitterfromn173_2 , buf_n173_splitterfromn173_1 , buf_n208_n211_1 , buf_n232_G2563_5 , buf_n232_G2563_4 , buf_n232_G2563_3 , buf_n232_G2563_2 , buf_n232_G2563_1 , buf_n233_n234_10 , buf_n233_n234_9 , buf_n233_n234_8 , buf_n233_n234_7 , buf_n233_n234_6 , buf_n233_n234_5 , buf_n233_n234_4 , buf_n233_n234_3 , buf_n233_n234_2 , buf_n233_n234_1 , buf_n236_n237_11 , buf_n236_n237_10 , buf_n236_n237_9 , buf_n236_n237_8 , buf_n236_n237_7 , buf_n236_n237_6 , buf_n236_n237_5 , buf_n236_n237_4 , buf_n236_n237_3 , buf_n236_n237_2 , buf_n236_n237_1 , buf_n237_G2565_1 , buf_n278_splitterfromn278_2 , buf_n278_splitterfromn278_1 , buf_n281_splitterfromn281_1 , buf_n282_n283_1 , buf_n283_G2577_4 , buf_n283_G2577_3 , buf_n283_G2577_2 , buf_n283_G2577_1 , buf_n287_splitterfromn287_4 , buf_n287_splitterfromn287_3 , buf_n287_splitterfromn287_2 , buf_n287_splitterfromn287_1 , buf_n298_G2580_8 , buf_n298_G2580_7 , buf_n298_G2580_6 , buf_n298_G2580_5 , buf_n298_G2580_4 , buf_n298_G2580_3 , buf_n298_G2580_2 , buf_n298_G2580_1 , buf_n299_n308_2 , buf_n299_n308_1 , buf_n310_n312_3 , buf_n310_n312_2 , buf_n310_n312_1 , buf_n314_n316_2 , buf_n314_n316_1 , buf_n320_n322_2 , buf_n320_n322_1 , buf_n324_n326_1 , buf_n329_n331_2 , buf_n329_n331_1 , buf_n335_n337_2 , buf_n335_n337_1 , buf_n339_n341_4 , buf_n339_n341_3 , buf_n339_n341_2 , buf_n339_n341_1 , buf_n352_n361_3 , buf_n352_n361_2 , buf_n352_n361_1 , buf_n386_n395_3 , buf_n386_n395_2 , buf_n386_n395_1 , buf_n398_n400_2 , buf_n398_n400_1 , buf_n404_n406_1 , buf_n410_n411_4 , buf_n410_n411_3 , buf_n410_n411_2 , buf_n410_n411_1 , buf_n420_n422_2 , buf_n420_n422_1 , buf_n428_splitterfromn428_3 , buf_n428_splitterfromn428_2 , buf_n428_splitterfromn428_1 , buf_n436_splitterfromn436_2 , buf_n436_splitterfromn436_1 , buf_n438_G2586_5 , buf_n438_G2586_4 , buf_n438_G2586_3 , buf_n438_G2586_2 , buf_n438_G2586_1 , buf_n445_splitterfromn445_4 , buf_n445_splitterfromn445_3 , buf_n445_splitterfromn445_2 , buf_n445_splitterfromn445_1 , buf_n447_splitterfromn447_2 , buf_n447_splitterfromn447_1 , buf_n452_n498_5 , buf_n452_n498_4 , buf_n452_n498_3 , buf_n452_n498_2 , buf_n452_n498_1 , buf_n454_n497_2 , buf_n454_n497_1 , buf_n455_n496_4 , buf_n455_n496_3 , buf_n455_n496_2 , buf_n455_n496_1 , buf_n517_n518_3 , buf_n517_n518_2 , buf_n517_n518_1 , buf_n522_n523_3 , buf_n522_n523_2 , buf_n522_n523_1 , buf_splitterfromG10_G2581_2 , buf_splitterfromG10_G2581_1 , buf_splitterfromG106_G2540_6 , buf_splitterfromG106_G2540_5 , buf_splitterfromG106_G2540_4 , buf_splitterfromG106_G2540_3 , buf_splitterfromG106_G2540_2 , buf_splitterfromG106_G2540_1 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_12 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_11 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_10 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_9 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_8 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_7 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_6 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_5 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_4 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_3 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_2 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_1 , buf_splitterfromG118_n282_1 , buf_splitterG123ton284n447_splitterG123ton276n447_1 , buf_splitterfromG125_n468_1 , buf_splitterfromG129_n456_2 , buf_splitterfromG129_n456_1 , buf_splitterfromG130_n480_2 , buf_splitterfromG130_n480_1 , buf_splitterG131ton368n487_n487_1 , buf_splitterfromG132_n455_1 , buf_splitterfromG133_n452_1 , buf_splitterG136ton500n469_splitterG136ton362n469_1 , buf_splitterG136ton362n469_n469_1 , buf_splitterG140ton327n457_n457_1 , buf_splitterG141ton158n481_n481_2 , buf_splitterG141ton158n481_n481_1 , buf_splitterG142ton332n488_n488_2 , buf_splitterG142ton332n488_n488_1 , buf_splitterfromG32_G2539_6 , buf_splitterfromG32_G2539_5 , buf_splitterfromG32_G2539_4 , buf_splitterfromG32_G2539_3 , buf_splitterfromG32_G2539_2 , buf_splitterfromG32_G2539_1 , buf_splitterfromG43_G2545_7 , buf_splitterfromG43_G2545_6 , buf_splitterfromG43_G2545_5 , buf_splitterfromG43_G2545_4 , buf_splitterfromG43_G2545_3 , buf_splitterfromG43_G2545_2 , buf_splitterfromG43_G2545_1 , buf_splitterfromG53_G2543_7 , buf_splitterfromG53_G2543_6 , buf_splitterfromG53_G2543_5 , buf_splitterfromG53_G2543_4 , buf_splitterfromG53_G2543_3 , buf_splitterfromG53_G2543_2 , buf_splitterfromG53_G2543_1 , buf_splitterfromG64_G2541_7 , buf_splitterfromG64_G2541_6 , buf_splitterfromG64_G2541_5 , buf_splitterfromG64_G2541_4 , buf_splitterfromG64_G2541_3 , buf_splitterfromG64_G2541_2 , buf_splitterfromG64_G2541_1 , buf_splitterfromG76_G2542_7 , buf_splitterfromG76_G2542_6 , buf_splitterfromG76_G2542_5 , buf_splitterfromG76_G2542_4 , buf_splitterfromG76_G2542_3 , buf_splitterfromG76_G2542_2 , buf_splitterfromG76_G2542_1 , buf_splitterfromG86_G2546_6 , buf_splitterfromG86_G2546_5 , buf_splitterfromG86_G2546_4 , buf_splitterfromG86_G2546_3 , buf_splitterfromG86_G2546_2 , buf_splitterfromG86_G2546_1 , buf_splitterfromG96_G2544_6 , buf_splitterfromG96_G2544_5 , buf_splitterfromG96_G2544_4 , buf_splitterfromG96_G2544_3 , buf_splitterfromG96_G2544_2 , buf_splitterfromG96_G2544_1 , buf_splittern164ton165G2551_G2551_4 , buf_splittern164ton165G2551_G2551_3 , buf_splittern164ton165G2551_G2551_2 , buf_splittern164ton165G2551_G2551_1 , buf_splittern176ton524G2556_G2556_1 , buf_splittern184ton345G2557_splittern184ton442G2557_2 , buf_splittern184ton345G2557_splittern184ton442G2557_1 , buf_splittern184ton442G2557_G2557_8 , buf_splittern184ton442G2557_G2557_7 , buf_splittern184ton442G2557_G2557_6 , buf_splittern184ton442G2557_G2557_5 , buf_splittern184ton442G2557_G2557_4 , buf_splittern184ton442G2557_G2557_3 , buf_splittern184ton442G2557_G2557_2 , buf_splittern184ton442G2557_G2557_1 , buf_splittern191ton330G2558_G2558_9 , buf_splittern191ton330G2558_G2558_8 , buf_splittern191ton330G2558_G2558_7 , buf_splittern191ton330G2558_G2558_6 , buf_splittern191ton330G2558_G2558_5 , buf_splittern191ton330G2558_G2558_4 , buf_splittern191ton330G2558_G2558_3 , buf_splittern191ton330G2558_G2558_2 , buf_splittern191ton330G2558_G2558_1 , buf_splittern198ton325G2559_G2559_10 , buf_splittern198ton325G2559_G2559_9 , buf_splittern198ton325G2559_G2559_8 , buf_splittern198ton325G2559_G2559_7 , buf_splittern198ton325G2559_G2559_6 , buf_splittern198ton325G2559_G2559_5 , buf_splittern198ton325G2559_G2559_4 , buf_splittern198ton325G2559_G2559_3 , buf_splittern198ton325G2559_G2559_2 , buf_splittern198ton325G2559_G2559_1 , buf_splittern207ton366G2569_splittern207ton486G2569_2 , buf_splittern207ton366G2569_splittern207ton486G2569_1 , buf_splittern207ton486G2569_splittern207toG2560G2569_6 , buf_splittern207ton486G2569_splittern207toG2560G2569_5 , buf_splittern207ton486G2569_splittern207toG2560G2569_4 , buf_splittern207ton486G2569_splittern207toG2560G2569_3 , buf_splittern207ton486G2569_splittern207toG2560G2569_2 , buf_splittern207ton486G2569_splittern207toG2560G2569_1 , buf_splittern215ton315G2568_splittern215ton479G2568_2 , buf_splittern215ton315G2568_splittern215ton479G2568_1 , buf_splittern215ton479G2568_splittern215ton280G2568_2 , buf_splittern215ton479G2568_splittern215ton280G2568_1 , buf_splittern215ton280G2568_splittern215toG2561G2568_3 , buf_splittern215ton280G2568_splittern215toG2561G2568_2 , buf_splittern215ton280G2568_splittern215toG2561G2568_1 , buf_splittern223ton321G2567_splittern223ton459G2567_3 , buf_splittern223ton321G2567_splittern223ton459G2567_2 , buf_splittern223ton321G2567_splittern223ton459G2567_1 , buf_splittern223ton277G2567_splittern223toG2562G2567_4 , buf_splittern223ton277G2567_splittern223toG2562G2567_3 , buf_splittern223ton277G2567_splittern223toG2562G2567_2 , buf_splittern223ton277G2567_splittern223toG2562G2567_1 , buf_splittern231ton311n232_splittern231ton284n232_2 , buf_splittern231ton311n232_splittern231ton284n232_1 , buf_splittern245ton336G2566_splittern245ton474G2566_2 , buf_splittern245ton336G2566_splittern245ton474G2566_1 , buf_splittern245ton474G2566_splittern245ton279G2566_1 , buf_splittern245ton279G2566_G2566_4 , buf_splittern245ton279G2566_G2566_3 , buf_splittern245ton279G2566_G2566_2 , buf_splittern245ton279G2566_G2566_1 , buf_splittern251ton421G2570_splittern251ton493G2570_4 , buf_splittern251ton421G2570_splittern251ton493G2570_3 , buf_splittern251ton421G2570_splittern251ton493G2570_2 , buf_splittern251ton421G2570_splittern251ton493G2570_1 , buf_splittern251ton493G2570_G2570_5 , buf_splittern251ton493G2570_G2570_4 , buf_splittern251ton493G2570_G2570_3 , buf_splittern251ton493G2570_G2570_2 , buf_splittern251ton493G2570_G2570_1 , buf_splittern259ton405G2571_splittern259ton454G2571_4 , buf_splittern259ton405G2571_splittern259ton454G2571_3 , buf_splittern259ton405G2571_splittern259ton454G2571_2 , buf_splittern259ton405G2571_splittern259ton454G2571_1 , buf_splittern259ton454G2571_G2571_5 , buf_splittern259ton454G2571_G2571_4 , buf_splittern259ton454G2571_G2571_3 , buf_splittern259ton454G2571_G2571_2 , buf_splittern259ton454G2571_G2571_1 , buf_splittern267ton399G2572_G2572_9 , buf_splittern267ton399G2572_G2572_8 , buf_splittern267ton399G2572_G2572_7 , buf_splittern267ton399G2572_G2572_6 , buf_splittern267ton399G2572_G2572_5 , buf_splittern267ton399G2572_G2572_4 , buf_splittern267ton399G2572_G2572_3 , buf_splittern267ton399G2572_G2572_2 , buf_splittern267ton399G2572_G2572_1 , buf_splittern275ton340n283_splittern275ton286n283_1 , buf_splitterfromn436_n446_2 , buf_splitterfromn436_n446_1 , buf_splitterfromn445_G2587_1 , buf_splittern453ton481n454_splittern453ton493n454_1 , buf_splittern503ton504n522_n522_2 , buf_splittern503ton504n522_n522_1 , buf_splitterfromn505_n519_1 , splitterfromG10 , splitterfromG106 , splitterG115ton163G2549 , splitterG115toG2531G2549 , splitterG117ton203n429 , splitterG117ton199n217 , splitterG117ton269n429 , splitterG117ton209n238 , splitterG117ton239n253 , splitterG117ton260n429 , splitterG117ton224n429 , splitterfromG118 , splitterfromG119 , splitterG12ton310n421 , splitterG12ton314n421 , splitterG12ton335n421 , splitterG12ton365n421 , splitterG12ton321n421 , splitterG12ton340n421 , splitterG120ton203n431 , splitterG120ton262n431 , splitterG120ton270n431 , splitterG120ton240n431 , splitterG121ton161n233 , splitterG122ton437n438 , splitterG122ton282n438 , splitterG123ton285n447 , splitterG123ton284n447 , splitterG123ton276n447 , splitterG123ton446n447 , splitterfromG124 , splitterfromG125 , splitterfromG126 , splitterfromG128 , splitterfromG129 , splitterfromG130 , splitterG131ton368n487 , splitterfromG132 , splitterfromG133 , splitterG134ton513n401 , splitterG134ton506n401 , splitterG135ton505n309 , splitterG135ton510n309 , splitterG136ton500n469 , splitterG136ton362n469 , splitterG137toG2536G2538 , splitterG138ton502n465 , splitterG138ton381n465 , splitterG139ton159n461 , splitterG139ton396n461 , splitterG140ton159n457 , splitterG140ton327n457 , splitterG141ton158n481 , splitterG142ton158n488 , splitterG142ton332n488 , splitterfromG143 , splitterfromG147 , splitterG23ton409n408 , splitterG23ton352n408 , splitterG23ton299n408 , splitterG23ton344n408 , splitterG23ton371n408 , splitterG23ton330n408 , splitterfromG32 , splitterfromG43 , splitterfromG53 , splitterfromG64 , splitterfromG76 , splitterG8ton451n486 , splitterG8ton479n486 , splitterfromG86 , splitterfromG96 , splittern164ton165G2551 , splitterfromn169 , splitterfromn172 , splitterfromn173 , splittern176ton234G2556 , splittern176ton524G2556 , splittern177ton178n391 , splittern177ton181n193 , splittern177ton195n391 , splittern177ton373n291 , splittern177ton185n188 , splittern177ton189n291 , splittern177ton292n391 , splittern177ton292n303 , splittern177ton304n356 , splittern177ton357n376 , splittern177ton387n391 , splittern184ton345G2557 , splittern184ton442G2557 , splittern191ton330G2558 , splittern198ton325G2559 , splittern203ton204n434 , splittern203ton205n220 , splittern203ton221n246 , splittern203ton264n434 , splittern203ton242n257 , splittern203ton272n434 , splittern207ton366G2569 , splittern207ton486G2569 , splittern207toG2560G2569 , splittern215ton315G2568 , splittern215ton479G2568 , splittern215ton280G2568 , splittern215toG2561G2568 , splittern223ton321G2567 , splittern223ton459G2567 , splittern223ton277G2567 , splittern223toG2562G2567 , splittern231ton311n232 , splittern231ton284n232 , splittern231ton471n232 , splitterfromn234 , splittern245ton336G2566 , splittern245ton474G2566 , splittern245ton279G2566 , splittern251ton421G2570 , splittern251ton493G2570 , splittern259ton405G2571 , splittern259ton454G2571 , splittern267ton399G2572 , splittern275ton340n283 , splittern275ton286n283 , splittern275ton467n283 , splittern275ton276n283 , splitterfromn278 , splitterfromn281 , splitterfromn287 , splittern294ton295n440 , splittern294ton408n440 , splittern306ton307n510 , splitterfromn309 , splitterfromn313 , splitterfromn317 , splitterfromn323 , splitterfromn327 , splitterfromn332 , splitterfromn338 , splitterfromn342 , splitterfromn347 , splitterfromn359 , splitterfromn361 , splitterfromn367 , splitterfromn378 , splitterfromn380 , splitterfromn396 , splitterfromn401 , splitterfromn407 , splitterfromn428 , splitterfromn436 , splitterfromn441 , splitterfromn445 , splitterfromn447 , splitterfromn448 , splitterfromn449 , splittern450ton460n469 , splittern450ton451n469 , splittern450ton456n469 , splittern451ton452n487 , splittern453ton481n454 , splittern453ton493n454 , splitterfromn459 , splitterfromn462 , splitterfromn466 , splitterfromn483 , splitterfromn490 , splittern499ton514n512 , splittern499ton503n512 , splitterfromn500 , splittern503ton504n522 , splitterfromn504 , splitterfromn505 , splitterfromn512 , splitterfromn514 , splitterfromn525 ;

PI_AQFP G1_( clk_1 , G1 );
PI_AQFP G10_( clk_1 , G10 );
PI_AQFP G100_( clk_1 , G100 );
PI_AQFP G101_( clk_1 , G101 );
PI_AQFP G102_( clk_1 , G102 );
PI_AQFP G103_( clk_1 , G103 );
PI_AQFP G105_( clk_1 , G105 );
PI_AQFP G106_( clk_1 , G106 );
PI_AQFP G107_( clk_1 , G107 );
PI_AQFP G108_( clk_1 , G108 );
PI_AQFP G109_( clk_1 , G109 );
PI_AQFP G11_( clk_1 , G11 );
PI_AQFP G110_( clk_1 , G110 );
PI_AQFP G111_( clk_1 , G111 );
PI_AQFP G112_( clk_1 , G112 );
PI_AQFP G113_( clk_1 , G113 );
PI_AQFP G114_( clk_1 , G114 );
PI_AQFP G115_( clk_1 , G115 );
PI_AQFP G116_( clk_1 , G116 );
PI_AQFP G117_( clk_1 , G117 );
PI_AQFP G118_( clk_1 , G118 );
PI_AQFP G119_( clk_1 , G119 );
PI_AQFP G12_( clk_1 , G12 );
PI_AQFP G120_( clk_1 , G120 );
PI_AQFP G121_( clk_1 , G121 );
PI_AQFP G122_( clk_1 , G122 );
PI_AQFP G123_( clk_1 , G123 );
PI_AQFP G124_( clk_1 , G124 );
PI_AQFP G125_( clk_1 , G125 );
PI_AQFP G126_( clk_1 , G126 );
PI_AQFP G127_( clk_1 , G127 );
PI_AQFP G128_( clk_1 , G128 );
PI_AQFP G129_( clk_1 , G129 );
PI_AQFP G13_( clk_1 , G13 );
PI_AQFP G130_( clk_1 , G130 );
PI_AQFP G131_( clk_1 , G131 );
PI_AQFP G132_( clk_1 , G132 );
PI_AQFP G133_( clk_1 , G133 );
PI_AQFP G134_( clk_1 , G134 );
PI_AQFP G135_( clk_1 , G135 );
PI_AQFP G136_( clk_1 , G136 );
PI_AQFP G137_( clk_1 , G137 );
PI_AQFP G138_( clk_1 , G138 );
PI_AQFP G139_( clk_1 , G139 );
PI_AQFP G14_( clk_1 , G14 );
PI_AQFP G140_( clk_1 , G140 );
PI_AQFP G141_( clk_1 , G141 );
PI_AQFP G142_( clk_1 , G142 );
PI_AQFP G143_( clk_1 , G143 );
PI_AQFP G144_( clk_1 , G144 );
PI_AQFP G145_( clk_1 , G145 );
PI_AQFP G146_( clk_1 , G146 );
PI_AQFP G147_( clk_1 , G147 );
PI_AQFP G148_( clk_1 , G148 );
PI_AQFP G149_( clk_1 , G149 );
PI_AQFP G15_( clk_1 , G15 );
PI_AQFP G150_( clk_1 , G150 );
PI_AQFP G151_( clk_1 , G151 );
PI_AQFP G152_( clk_1 , G152 );
PI_AQFP G153_( clk_1 , G153 );
PI_AQFP G154_( clk_1 , G154 );
PI_AQFP G155_( clk_1 , G155 );
PI_AQFP G156_( clk_1 , G156 );
PI_AQFP G157_( clk_1 , G157 );
PI_AQFP G16_( clk_1 , G16 );
PI_AQFP G17_( clk_1 , G17 );
PI_AQFP G18_( clk_1 , G18 );
PI_AQFP G19_( clk_1 , G19 );
PI_AQFP G2_( clk_1 , G2 );
PI_AQFP G20_( clk_1 , G20 );
PI_AQFP G21_( clk_1 , G21 );
PI_AQFP G22_( clk_1 , G22 );
PI_AQFP G23_( clk_1 , G23 );
PI_AQFP G24_( clk_1 , G24 );
PI_AQFP G25_( clk_1 , G25 );
PI_AQFP G26_( clk_1 , G26 );
PI_AQFP G27_( clk_1 , G27 );
PI_AQFP G28_( clk_1 , G28 );
PI_AQFP G29_( clk_1 , G29 );
PI_AQFP G3_( clk_1 , G3 );
PI_AQFP G30_( clk_1 , G30 );
PI_AQFP G31_( clk_1 , G31 );
PI_AQFP G32_( clk_1 , G32 );
PI_AQFP G33_( clk_1 , G33 );
PI_AQFP G34_( clk_1 , G34 );
PI_AQFP G35_( clk_1 , G35 );
PI_AQFP G36_( clk_1 , G36 );
PI_AQFP G37_( clk_1 , G37 );
PI_AQFP G38_( clk_1 , G38 );
PI_AQFP G39_( clk_1 , G39 );
PI_AQFP G4_( clk_1 , G4 );
PI_AQFP G40_( clk_1 , G40 );
PI_AQFP G41_( clk_1 , G41 );
PI_AQFP G42_( clk_1 , G42 );
PI_AQFP G43_( clk_1 , G43 );
PI_AQFP G44_( clk_1 , G44 );
PI_AQFP G45_( clk_1 , G45 );
PI_AQFP G46_( clk_1 , G46 );
PI_AQFP G47_( clk_1 , G47 );
PI_AQFP G48_( clk_1 , G48 );
PI_AQFP G49_( clk_1 , G49 );
PI_AQFP G5_( clk_1 , G5 );
PI_AQFP G50_( clk_1 , G50 );
PI_AQFP G51_( clk_1 , G51 );
PI_AQFP G52_( clk_1 , G52 );
PI_AQFP G53_( clk_1 , G53 );
PI_AQFP G54_( clk_1 , G54 );
PI_AQFP G55_( clk_1 , G55 );
PI_AQFP G56_( clk_1 , G56 );
PI_AQFP G57_( clk_1 , G57 );
PI_AQFP G58_( clk_1 , G58 );
PI_AQFP G59_( clk_1 , G59 );
PI_AQFP G6_( clk_1 , G6 );
PI_AQFP G60_( clk_1 , G60 );
PI_AQFP G61_( clk_1 , G61 );
PI_AQFP G62_( clk_1 , G62 );
PI_AQFP G63_( clk_1 , G63 );
PI_AQFP G64_( clk_1 , G64 );
PI_AQFP G65_( clk_1 , G65 );
PI_AQFP G66_( clk_1 , G66 );
PI_AQFP G67_( clk_1 , G67 );
PI_AQFP G68_( clk_1 , G68 );
PI_AQFP G69_( clk_1 , G69 );
PI_AQFP G7_( clk_1 , G7 );
PI_AQFP G70_( clk_1 , G70 );
PI_AQFP G71_( clk_1 , G71 );
PI_AQFP G72_( clk_1 , G72 );
PI_AQFP G73_( clk_1 , G73 );
PI_AQFP G74_( clk_1 , G74 );
PI_AQFP G75_( clk_1 , G75 );
PI_AQFP G76_( clk_1 , G76 );
PI_AQFP G77_( clk_1 , G77 );
PI_AQFP G78_( clk_1 , G78 );
PI_AQFP G79_( clk_1 , G79 );
PI_AQFP G8_( clk_1 , G8 );
PI_AQFP G80_( clk_1 , G80 );
PI_AQFP G81_( clk_1 , G81 );
PI_AQFP G82_( clk_1 , G82 );
PI_AQFP G83_( clk_1 , G83 );
PI_AQFP G84_( clk_1 , G84 );
PI_AQFP G85_( clk_1 , G85 );
PI_AQFP G86_( clk_1 , G86 );
PI_AQFP G87_( clk_1 , G87 );
PI_AQFP G88_( clk_1 , G88 );
PI_AQFP G89_( clk_1 , G89 );
PI_AQFP G9_( clk_1 , G9 );
PI_AQFP G90_( clk_1 , G90 );
PI_AQFP G91_( clk_1 , G91 );
PI_AQFP G92_( clk_1 , G92 );
PI_AQFP G93_( clk_1 , G93 );
PI_AQFP G94_( clk_1 , G94 );
PI_AQFP G95_( clk_1 , G95 );
PI_AQFP G96_( clk_1 , G96 );
PI_AQFP G97_( clk_1 , G97 );
PI_AQFP G98_( clk_1 , G98 );
PI_AQFP G99_( clk_1 , G99 );
or_AQFP n158_( clk_3 , splitterG141ton158n481 , splitterG142ton158n488 , 0 , 0 , n158 );
or_AQFP n159_( clk_3 , splitterG139ton159n461 , splitterG140ton159n457 , 0 , 0 , n159 );
or_AQFP n160_( clk_5 , n158 , n159 , 0 , 0 , n160 );
or_AQFP n161_( clk_3 , splitterG121ton161n233 , G2 , 0 , 0 , n161 );
or_AQFP n162_( clk_4 , buf_G11_n162_1 , n161 , 0 , 0 , n162 );
and_AQFP n163_( clk_4 , splitterG115ton163G2549 , buf_G74_n163_1 , 0 , 1 , n163 );
or_AQFP n164_( clk_3 , splitterG121ton161n233 , G7 , 0 , 0 , n164 );
or_AQFP n165_( clk_6 , splitterfromG119 , splittern164ton165G2551 , 0 , 0 , n165 );
or_AQFP n166_( clk_6 , splitterfromG147 , splittern164ton165G2551 , 0 , 0 , n166 );
and_AQFP n167_( clk_1 , splitterfromG53 , splitterfromG96 , 0 , 1 , n167 );
or_AQFP n168_( clk_1 , splitterfromG43 , splitterfromG86 , 0 , 0 , n168 );
and_AQFP n169_( clk_3 , n167 , n168 , 0 , 1 , n169 );
and_AQFP n170_( clk_2 , splitterfromG106 , splitterfromG32 , 1 , 0 , n170 );
or_AQFP n171_( clk_1 , splitterfromG64 , splitterfromG76 , 0 , 0 , n171 );
and_AQFP n172_( clk_3 , n170 , n171 , 0 , 1 , n172 );
or_AQFP n173_( clk_7 , splitterfromn169 , splitterfromn172 , 0 , 0 , n173 );
and_AQFP n174_( clk_6 , splitterfromG147 , splitterfromn172 , 0 , 1 , n174 );
and_AQFP n175_( clk_6 , splitterfromG119 , splitterfromn169 , 0 , 1 , n175 );
or_AQFP n176_( clk_7 , n174 , n175 , 0 , 0 , n176 );
or_AQFP n177_( clk_2 , G145 , G146 , 0 , 0 , n177 );
and_AQFP n178_( clk_4 , buf_G109_n178_1 , splittern177ton178n391 , 0 , 1 , n178 );
and_AQFP n179_( clk_4 , buf_G79_n179_1 , splittern177ton178n391 , 0 , 1 , n179 );
or_AQFP n180_( clk_5 , n178 , n179 , 0 , 0 , n180 );
and_AQFP n181_( clk_5 , buf_G89_n181_1 , splittern177ton181n193 , 0 , 1 , n181 );
and_AQFP n182_( clk_5 , buf_G99_n182_1 , splittern177ton181n193 , 0 , 1 , n182 );
or_AQFP n183_( clk_6 , n181 , n182 , 0 , 0 , n183 );
or_AQFP n184_( clk_7 , n180 , n183 , 0 , 0 , n184 );
or_AQFP n185_( clk_7 , buf_G108_n185_1 , splittern177ton185n188 , 0 , 0 , n185 );
and_AQFP n186_( clk_7 , buf_G98_n186_1 , splittern177ton185n188 , 0 , 1 , n186 );
and_AQFP n187_( clk_8 , n185 , n186 , 0 , 1 , n187 );
and_AQFP n188_( clk_7 , buf_G88_n188_1 , splittern177ton185n188 , 0 , 1 , n188 );
and_AQFP n189_( clk_7 , buf_G78_n189_1 , splittern177ton189n291 , 0 , 1 , n189 );
or_AQFP n190_( clk_8 , n188 , n189 , 0 , 0 , n190 );
and_AQFP n191_( clk_1 , n187 , n190 , 0 , 1 , n191 );
or_AQFP n192_( clk_5 , buf_G80_n192_1 , splittern177ton181n193 , 0 , 0 , n192 );
and_AQFP n193_( clk_5 , buf_G90_n193_1 , splittern177ton181n193 , 0 , 1 , n193 );
and_AQFP n194_( clk_6 , n192 , n193 , 0 , 1 , n194 );
and_AQFP n195_( clk_5 , buf_G100_n195_1 , splittern177ton195n391 , 0 , 1 , n195 );
and_AQFP n196_( clk_5 , buf_G110_n196_1 , splittern177ton195n391 , 0 , 1 , n196 );
or_AQFP n197_( clk_6 , n195 , n196 , 0 , 0 , n197 );
and_AQFP n198_( clk_7 , n194 , n197 , 0 , 1 , n198 );
and_AQFP n199_( clk_4 , splitterG117ton199n217 , buf_G36_n199_1 , 0 , 1 , n199 );
and_AQFP n200_( clk_4 , splitterG117ton199n217 , buf_G68_n200_1 , 0 , 1 , n200 );
or_AQFP n201_( clk_5 , splitterG120ton262n431 , n200 , 0 , 0 , n201 );
and_AQFP n202_( clk_6 , n199 , n201 , 0 , 1 , n202 );
or_AQFP n203_( clk_3 , splitterG117ton203n429 , splitterG120ton203n431 , 0 , 0 , n203 );
and_AQFP n204_( clk_5 , buf_G46_n204_1 , splittern203ton204n434 , 0 , 1 , n204 );
and_AQFP n205_( clk_6 , buf_G57_n205_1 , splittern203ton205n220 , 0 , 1 , n205 );
or_AQFP n206_( clk_7 , n204 , n205 , 0 , 0 , n206 );
and_AQFP n207_( clk_8 , n202 , n206 , 0 , 1 , n207 );
and_AQFP n208_( clk_4 , splitterG117ton199n217 , buf_G37_n208_1 , 0 , 1 , n208 );
and_AQFP n209_( clk_5 , splitterG117ton209n238 , buf_G69_n209_1 , 0 , 1 , n209 );
or_AQFP n210_( clk_6 , splitterG120ton270n431 , n209 , 0 , 0 , n210 );
and_AQFP n211_( clk_7 , buf_n208_n211_1 , n210 , 0 , 1 , n211 );
and_AQFP n212_( clk_6 , buf_G47_n212_1 , splittern203ton205n220 , 0 , 1 , n212 );
and_AQFP n213_( clk_6 , buf_G58_n213_1 , splittern203ton205n220 , 0 , 1 , n213 );
or_AQFP n214_( clk_7 , n212 , n213 , 0 , 0 , n214 );
and_AQFP n215_( clk_8 , n211 , n214 , 0 , 1 , n215 );
and_AQFP n216_( clk_5 , splitterG117ton209n238 , buf_G38_n216_1 , 0 , 1 , n216 );
and_AQFP n217_( clk_4 , splitterG117ton199n217 , buf_G70_n217_1 , 0 , 1 , n217 );
or_AQFP n218_( clk_5 , splitterG120ton262n431 , n217 , 0 , 0 , n218 );
and_AQFP n219_( clk_6 , n216 , n218 , 0 , 1 , n219 );
and_AQFP n220_( clk_6 , buf_G48_n220_1 , splittern203ton205n220 , 0 , 1 , n220 );
and_AQFP n221_( clk_6 , buf_G59_n221_1 , splittern203ton221n246 , 0 , 1 , n221 );
or_AQFP n222_( clk_7 , n220 , n221 , 0 , 0 , n222 );
and_AQFP n223_( clk_8 , n219 , n222 , 0 , 1 , n223 );
and_AQFP n224_( clk_6 , splitterG117ton224n429 , buf_G31_n224_1 , 0 , 1 , n224 );
and_AQFP n225_( clk_5 , splitterG117ton209n238 , buf_G63_n225_1 , 0 , 1 , n225 );
or_AQFP n226_( clk_6 , splitterG120ton270n431 , n225 , 0 , 0 , n226 );
and_AQFP n227_( clk_7 , n224 , n226 , 0 , 1 , n227 );
and_AQFP n228_( clk_6 , buf_G42_n228_1 , splittern203ton221n246 , 0 , 1 , n228 );
and_AQFP n229_( clk_6 , buf_G52_n229_1 , splittern203ton221n246 , 0 , 1 , n229 );
or_AQFP n230_( clk_7 , n228 , n229 , 0 , 0 , n230 );
and_AQFP n231_( clk_8 , n227 , n230 , 0 , 1 , n231 );
or_AQFP n232_( clk_2 , splitterG122ton282n438 , splittern231ton471n232 , 0 , 0 , n232 );
or_AQFP n233_( clk_4 , buf_G116_n233_1 , splitterG121ton161n233 , 0 , 0 , n233 );
or_AQFP n234_( clk_1 , splittern176ton234G2556 , buf_n233_n234_1 , 0 , 0 , n234 );
or_AQFP n235_( clk_4 , buf_G28_n235_1 , splitterfromn234 , 0 , 0 , n235 );
and_AQFP n236_( clk_3 , G1 , G3 , 0 , 1 , n236 );
or_AQFP n237_( clk_3 , splitterfromn234 , buf_n236_n237_1 , 0 , 0 , n237 );
or_AQFP n238_( clk_5 , splitterG117ton209n238 , buf_G39_n238_1 , 0 , 0 , n238 );
and_AQFP n239_( clk_5 , splitterG117ton239n253 , buf_G71_n239_1 , 0 , 1 , n239 );
or_AQFP n240_( clk_6 , splitterG120ton240n431 , n239 , 0 , 0 , n240 );
and_AQFP n241_( clk_7 , n238 , n240 , 0 , 1 , n241 );
and_AQFP n242_( clk_7 , buf_G49_n242_1 , splittern203ton242n257 , 0 , 1 , n242 );
and_AQFP n243_( clk_7 , buf_G60_n243_1 , splittern203ton242n257 , 0 , 1 , n243 );
or_AQFP n244_( clk_8 , n242 , n243 , 0 , 0 , n244 );
or_AQFP n245_( clk_1 , n241 , n244 , 0 , 0 , n245 );
and_AQFP n246_( clk_6 , buf_G56_n246_1 , splittern203ton221n246 , 0 , 1 , n246 );
or_AQFP n247_( clk_6 , splitterG117ton224n429 , buf_G35_n247_1 , 0 , 0 , n247 );
and_AQFP n248_( clk_5 , splitterG117ton239n253 , buf_G67_n248_1 , 0 , 1 , n248 );
or_AQFP n249_( clk_6 , splitterG120ton240n431 , n248 , 0 , 0 , n249 );
and_AQFP n250_( clk_7 , n247 , n249 , 0 , 1 , n250 );
and_AQFP n251_( clk_8 , n246 , n250 , 0 , 1 , n251 );
and_AQFP n252_( clk_5 , splitterG117ton239n253 , buf_G34_n252_1 , 0 , 1 , n252 );
and_AQFP n253_( clk_5 , splitterG117ton239n253 , buf_G66_n253_1 , 0 , 1 , n253 );
or_AQFP n254_( clk_6 , splitterG120ton240n431 , n253 , 0 , 0 , n254 );
and_AQFP n255_( clk_7 , n252 , n254 , 0 , 1 , n255 );
and_AQFP n256_( clk_7 , buf_G45_n256_1 , splittern203ton242n257 , 0 , 1 , n256 );
and_AQFP n257_( clk_7 , buf_G55_n257_1 , splittern203ton242n257 , 0 , 1 , n257 );
or_AQFP n258_( clk_8 , n256 , n257 , 0 , 0 , n258 );
and_AQFP n259_( clk_1 , n255 , n258 , 0 , 1 , n259 );
and_AQFP n260_( clk_5 , splitterG117ton260n429 , buf_G33_n260_1 , 0 , 1 , n260 );
and_AQFP n261_( clk_3 , splitterG117ton203n429 , G65 , 0 , 1 , n261 );
or_AQFP n262_( clk_4 , splitterG120ton262n431 , n261 , 0 , 0 , n262 );
and_AQFP n263_( clk_6 , n260 , n262 , 0 , 1 , n263 );
and_AQFP n264_( clk_6 , buf_G44_n264_1 , splittern203ton264n434 , 0 , 1 , n264 );
and_AQFP n265_( clk_6 , buf_G54_n265_1 , splittern203ton264n434 , 0 , 1 , n265 );
or_AQFP n266_( clk_7 , n264 , n265 , 0 , 0 , n266 );
and_AQFP n267_( clk_8 , n263 , n266 , 0 , 1 , n267 );
and_AQFP n268_( clk_5 , splitterG117ton260n429 , buf_G40_n268_1 , 0 , 1 , n268 );
and_AQFP n269_( clk_4 , splitterG117ton269n429 , buf_G72_n269_1 , 0 , 1 , n269 );
or_AQFP n270_( clk_5 , splitterG120ton270n431 , n269 , 0 , 0 , n270 );
and_AQFP n271_( clk_7 , n268 , n270 , 0 , 1 , n271 );
and_AQFP n272_( clk_7 , buf_G50_n272_1 , splittern203ton272n434 , 0 , 1 , n272 );
and_AQFP n273_( clk_7 , buf_G61_n273_1 , splittern203ton272n434 , 0 , 1 , n273 );
or_AQFP n274_( clk_8 , n272 , n273 , 0 , 0 , n274 );
and_AQFP n275_( clk_1 , n271 , n274 , 0 , 1 , n275 );
or_AQFP n276_( clk_4 , splitterG123ton276n447 , splittern275ton276n283 , 0 , 0 , n276 );
and_AQFP n277_( clk_4 , splitterG123ton276n447 , splittern223ton277G2567 , 0 , 1 , n277 );
and_AQFP n278_( clk_6 , n276 , n277 , 0 , 1 , n278 );
or_AQFP n279_( clk_6 , splitterG123ton446n447 , splittern245ton279G2566 , 0 , 0 , n279 );
and_AQFP n280_( clk_6 , splitterG123ton446n447 , splittern215ton280G2568 , 1 , 0 , n280 );
and_AQFP n281_( clk_8 , n279 , n280 , 0 , 1 , n281 );
and_AQFP n282_( clk_1 , buf_splitterfromG118_n282_1 , splitterG122ton282n438 , 0 , 1 , n282 );
or_AQFP n283_( clk_4 , splittern275ton276n283 , buf_n282_n283_1 , 0 , 0 , n283 );
and_AQFP n284_( clk_8 , splitterG123ton284n447 , splittern231ton284n232 , 0 , 1 , n284 );
or_AQFP n285_( clk_6 , splitterfromG118 , splitterG123ton285n447 , 0 , 0 , n285 );
and_AQFP n286_( clk_8 , splittern275ton286n283 , n285 , 0 , 1 , n286 );
or_AQFP n287_( clk_2 , n284 , n286 , 0 , 0 , n287 );
and_AQFP n288_( clk_7 , buf_G77_n288_1 , splittern177ton189n291 , 0 , 1 , n288 );
and_AQFP n289_( clk_7 , buf_G97_n289_1 , splittern177ton189n291 , 0 , 1 , n289 );
and_AQFP n290_( clk_8 , n288 , n289 , 0 , 1 , n290 );
and_AQFP n291_( clk_7 , buf_G107_n291_1 , splittern177ton189n291 , 0 , 1 , n291 );
and_AQFP n292_( clk_7 , buf_G87_n292_1 , splittern177ton292n303 , 0 , 1 , n292 );
or_AQFP n293_( clk_8 , n291 , n292 , 0 , 0 , n293 );
and_AQFP n294_( clk_1 , n290 , n293 , 0 , 1 , n294 );
or_AQFP n295_( clk_3 , splitterfromG143 , splittern294ton295n440 , 0 , 0 , n295 );
and_AQFP n296_( clk_3 , splitterfromG143 , splittern294ton295n440 , 0 , 1 , n296 );
and_AQFP n297_( clk_4 , n295 , n296 , 0 , 1 , n297 );
or_AQFP n298_( clk_5 , buf_G144_n298_1 , n297 , 0 , 0 , n298 );
and_AQFP n299_( clk_7 , buf_G19_n299_1 , splitterG23ton299n408 , 1 , 0 , n299 );
and_AQFP n300_( clk_7 , buf_G75_n300_1 , splittern177ton292n303 , 0 , 1 , n300 );
and_AQFP n301_( clk_7 , buf_G85_n301_1 , splittern177ton292n303 , 0 , 1 , n301 );
and_AQFP n302_( clk_8 , n300 , n301 , 0 , 1 , n302 );
and_AQFP n303_( clk_7 , buf_G95_n303_1 , splittern177ton292n303 , 0 , 1 , n303 );
and_AQFP n304_( clk_7 , buf_G105_n304_1 , splittern177ton304n356 , 0 , 1 , n304 );
or_AQFP n305_( clk_8 , n303 , n304 , 0 , 0 , n305 );
and_AQFP n306_( clk_1 , n302 , n305 , 0 , 1 , n306 );
and_AQFP n307_( clk_3 , splitterG23ton371n408 , splittern306ton307n510 , 0 , 1 , n307 );
and_AQFP n308_( clk_4 , buf_n299_n308_1 , n307 , 0 , 1 , n308 );
and_AQFP n309_( clk_5 , splitterG135ton510n309 , n308 , 0 , 1 , n309 );
and_AQFP n310_( clk_3 , splitterG12ton310n421 , G13 , 0 , 1 , n310 );
and_AQFP n311_( clk_2 , splitterG12ton365n421 , splittern231ton311n232 , 0 , 1 , n311 );
and_AQFP n312_( clk_3 , buf_n310_n312_1 , n311 , 0 , 1 , n312 );
and_AQFP n313_( clk_5 , splitterfromG125 , n312 , 0 , 1 , n313 );
and_AQFP n314_( clk_5 , splitterG12ton314n421 , buf_G15_n314_1 , 0 , 1 , n314 );
and_AQFP n315_( clk_2 , splitterG12ton365n421 , splittern215ton315G2568 , 1 , 0 , n315 );
and_AQFP n316_( clk_3 , buf_n314_n316_1 , n315 , 0 , 1 , n316 );
and_AQFP n317_( clk_4 , splitterfromG130 , n316 , 0 , 1 , n317 );
or_AQFP n318_( clk_7 , splitterfromn313 , splitterfromn317 , 0 , 0 , n318 );
or_AQFP n319_( clk_1 , splitterfromn309 , n318 , 0 , 0 , n319 );
and_AQFP n320_( clk_5 , splitterG12ton314n421 , buf_G5_n320_1 , 0 , 1 , n320 );
and_AQFP n321_( clk_2 , splitterG12ton321n421 , splittern223ton321G2567 , 0 , 1 , n321 );
and_AQFP n322_( clk_3 , buf_n320_n322_1 , n321 , 0 , 1 , n322 );
and_AQFP n323_( clk_4 , splitterfromG129 , n322 , 0 , 1 , n323 );
and_AQFP n324_( clk_6 , buf_G21_n324_1 , splitterG23ton299n408 , 1 , 0 , n324 );
and_AQFP n325_( clk_1 , splitterG23ton344n408 , splittern198ton325G2559 , 0 , 1 , n325 );
and_AQFP n326_( clk_2 , buf_n324_n326_1 , n325 , 0 , 1 , n326 );
and_AQFP n327_( clk_4 , splitterG140ton327n457 , n326 , 0 , 1 , n327 );
or_AQFP n328_( clk_7 , splitterfromn323 , splitterfromn327 , 0 , 0 , n328 );
and_AQFP n329_( clk_6 , splitterG23ton299n408 , buf_G27_n329_1 , 0 , 1 , n329 );
and_AQFP n330_( clk_3 , splitterG23ton330n408 , splittern191ton330G2558 , 0 , 1 , n330 );
and_AQFP n331_( clk_4 , buf_n329_n331_1 , n330 , 0 , 1 , n331 );
and_AQFP n332_( clk_5 , splitterG142ton332n488 , n331 , 0 , 1 , n332 );
or_AQFP n333_( clk_8 , splitterfromn309 , splitterfromn332 , 0 , 0 , n333 );
or_AQFP n334_( clk_1 , n328 , n333 , 0 , 0 , n334 );
and_AQFP n335_( clk_7 , splitterG12ton335n421 , buf_G14_n335_1 , 0 , 1 , n335 );
and_AQFP n336_( clk_3 , splitterG12ton321n421 , splittern245ton336G2566 , 1 , 0 , n336 );
and_AQFP n337_( clk_4 , buf_n335_n337_1 , n336 , 0 , 1 , n337 );
and_AQFP n338_( clk_5 , splitterfromG128 , n337 , 0 , 1 , n338 );
and_AQFP n339_( clk_3 , splitterG12ton310n421 , G4 , 0 , 1 , n339 );
and_AQFP n340_( clk_3 , splitterG12ton340n421 , splittern275ton340n283 , 0 , 1 , n340 );
and_AQFP n341_( clk_4 , buf_n339_n341_1 , n340 , 0 , 1 , n341 );
and_AQFP n342_( clk_5 , splitterfromG126 , n341 , 0 , 1 , n342 );
or_AQFP n343_( clk_7 , splitterfromn338 , splitterfromn342 , 0 , 0 , n343 );
and_AQFP n344_( clk_8 , splitterG23ton344n408 , buf_G26_n344_1 , 0 , 1 , n344 );
and_AQFP n345_( clk_1 , splitterG23ton344n408 , splittern184ton345G2557 , 0 , 1 , n345 );
and_AQFP n346_( clk_2 , n344 , n345 , 0 , 1 , n346 );
and_AQFP n347_( clk_3 , splitterG141ton158n481 , n346 , 0 , 1 , n347 );
or_AQFP n348_( clk_6 , splitterfromn327 , splitterfromn347 , 0 , 0 , n348 );
or_AQFP n349_( clk_8 , n343 , n348 , 0 , 0 , n349 );
or_AQFP n350_( clk_2 , n334 , n349 , 0 , 0 , n350 );
or_AQFP n351_( clk_3 , n319 , n350 , 0 , 0 , n351 );
and_AQFP n352_( clk_4 , splitterG23ton352n408 , buf_G24_n352_1 , 0 , 1 , n352 );
and_AQFP n353_( clk_7 , buf_G93_n353_1 , splittern177ton304n356 , 0 , 1 , n353 );
and_AQFP n354_( clk_7 , buf_G103_n354_1 , splittern177ton304n356 , 0 , 1 , n354 );
and_AQFP n355_( clk_8 , n353 , n354 , 0 , 1 , n355 );
and_AQFP n356_( clk_7 , buf_G113_n356_1 , splittern177ton304n356 , 0 , 1 , n356 );
and_AQFP n357_( clk_7 , buf_G83_n357_1 , splittern177ton357n376 , 0 , 1 , n357 );
or_AQFP n358_( clk_8 , n356 , n357 , 0 , 0 , n358 );
and_AQFP n359_( clk_1 , n355 , n358 , 0 , 1 , n359 );
and_AQFP n360_( clk_3 , splitterG23ton330n408 , splitterfromn359 , 0 , 1 , n360 );
and_AQFP n361_( clk_4 , buf_n352_n361_1 , n360 , 0 , 1 , n361 );
or_AQFP n362_( clk_6 , splitterG136ton362n469 , splitterfromn361 , 0 , 0 , n362 );
and_AQFP n363_( clk_6 , splitterG136ton362n469 , splitterfromn361 , 0 , 1 , n363 );
and_AQFP n364_( clk_7 , n362 , n363 , 0 , 1 , n364 );
and_AQFP n365_( clk_1 , splitterG12ton365n421 , buf_G16_n365_1 , 0 , 1 , n365 );
and_AQFP n366_( clk_2 , splitterG12ton321n421 , splittern207ton366G2569 , 0 , 1 , n366 );
and_AQFP n367_( clk_3 , n365 , n366 , 0 , 1 , n367 );
or_AQFP n368_( clk_5 , splitterG131ton368n487 , splitterfromn367 , 0 , 0 , n368 );
and_AQFP n369_( clk_5 , splitterG131ton368n487 , splitterfromn367 , 0 , 1 , n369 );
and_AQFP n370_( clk_6 , n368 , n369 , 0 , 1 , n370 );
and_AQFP n371_( clk_2 , buf_G20_n371_1 , splitterG23ton371n408 , 1 , 0 , n371 );
and_AQFP n372_( clk_7 , buf_G82_n372_1 , splittern177ton357n376 , 0 , 1 , n372 );
and_AQFP n373_( clk_6 , buf_G102_n373_1 , splittern177ton373n291 , 0 , 1 , n373 );
and_AQFP n374_( clk_8 , n372 , n373 , 0 , 1 , n374 );
and_AQFP n375_( clk_7 , buf_G112_n375_1 , splittern177ton357n376 , 0 , 1 , n375 );
and_AQFP n376_( clk_7 , buf_G92_n376_1 , splittern177ton357n376 , 0 , 1 , n376 );
or_AQFP n377_( clk_8 , n375 , n376 , 0 , 0 , n377 );
and_AQFP n378_( clk_1 , n374 , n377 , 0 , 1 , n378 );
and_AQFP n379_( clk_3 , splitterG23ton330n408 , splitterfromn378 , 0 , 1 , n379 );
and_AQFP n380_( clk_4 , n371 , n379 , 0 , 1 , n380 );
or_AQFP n381_( clk_6 , splitterG138ton381n465 , splitterfromn380 , 0 , 0 , n381 );
and_AQFP n382_( clk_6 , splitterG138ton381n465 , splitterfromn380 , 0 , 1 , n382 );
and_AQFP n383_( clk_7 , n381 , n382 , 0 , 1 , n383 );
or_AQFP n384_( clk_8 , n370 , n383 , 0 , 0 , n384 );
or_AQFP n385_( clk_1 , n364 , n384 , 0 , 0 , n385 );
and_AQFP n386_( clk_4 , splitterG23ton352n408 , buf_G25_n386_1 , 0 , 1 , n386 );
and_AQFP n387_( clk_7 , buf_G81_n387_1 , splittern177ton387n391 , 0 , 1 , n387 );
and_AQFP n388_( clk_7 , buf_G101_n388_1 , splittern177ton387n391 , 0 , 1 , n388 );
and_AQFP n389_( clk_8 , n387 , n388 , 0 , 1 , n389 );
and_AQFP n390_( clk_7 , buf_G111_n390_1 , splittern177ton387n391 , 0 , 1 , n390 );
and_AQFP n391_( clk_7 , buf_G91_n391_1 , splittern177ton387n391 , 0 , 1 , n391 );
or_AQFP n392_( clk_8 , n390 , n391 , 0 , 0 , n392 );
and_AQFP n393_( clk_1 , n389 , n392 , 0 , 1 , n393 );
and_AQFP n394_( clk_2 , splitterG23ton371n408 , n393 , 0 , 1 , n394 );
and_AQFP n395_( clk_3 , buf_n386_n395_1 , n394 , 0 , 1 , n395 );
and_AQFP n396_( clk_4 , splitterG139ton396n461 , n395 , 0 , 1 , n396 );
or_AQFP n397_( clk_6 , splitterfromn317 , splitterfromn396 , 0 , 0 , n397 );
and_AQFP n398_( clk_6 , splitterG12ton314n421 , buf_G18_n398_1 , 0 , 1 , n398 );
and_AQFP n399_( clk_3 , splitterG12ton340n421 , splittern267ton399G2572 , 0 , 1 , n399 );
and_AQFP n400_( clk_4 , buf_n398_n400_1 , n399 , 0 , 1 , n400 );
and_AQFP n401_( clk_5 , splitterG134ton506n401 , n400 , 0 , 1 , n401 );
or_AQFP n402_( clk_7 , splitterfromn342 , splitterfromn401 , 0 , 0 , n402 );
or_AQFP n403_( clk_8 , n397 , n402 , 0 , 0 , n403 );
and_AQFP n404_( clk_8 , splitterG12ton335n421 , buf_G6_n404_1 , 0 , 1 , n404 );
and_AQFP n405_( clk_3 , splitterG12ton340n421 , splittern259ton405G2571 , 0 , 1 , n405 );
and_AQFP n406_( clk_4 , buf_n404_n406_1 , n405 , 0 , 1 , n406 );
and_AQFP n407_( clk_5 , splitterfromG133 , n406 , 0 , 1 , n407 );
and_AQFP n408_( clk_4 , splitterG23ton330n408 , splittern294ton408n440 , 0 , 1 , n408 );
and_AQFP n409_( clk_3 , G22 , splitterG23ton409n408 , 1 , 0 , n409 );
or_AQFP n410_( clk_4 , buf_G9_n410_1 , n409 , 0 , 0 , n410 );
or_AQFP n411_( clk_5 , n408 , buf_n410_n411_1 , 0 , 0 , n411 );
or_AQFP n412_( clk_7 , splitterfromn407 , n411 , 0 , 0 , n412 );
or_AQFP n413_( clk_7 , splitterfromn332 , splitterfromn407 , 0 , 0 , n413 );
or_AQFP n414_( clk_8 , n412 , n413 , 0 , 0 , n414 );
or_AQFP n415_( clk_1 , n403 , n414 , 0 , 0 , n415 );
or_AQFP n416_( clk_6 , splitterfromn323 , splitterfromn347 , 0 , 0 , n416 );
or_AQFP n417_( clk_7 , splitterfromn313 , splitterfromn338 , 0 , 0 , n417 );
or_AQFP n418_( clk_8 , n416 , n417 , 0 , 0 , n418 );
or_AQFP n419_( clk_7 , splitterfromn396 , splitterfromn401 , 0 , 0 , n419 );
and_AQFP n420_( clk_7 , splitterG12ton335n421 , buf_G17_n420_1 , 0 , 1 , n420 );
and_AQFP n421_( clk_3 , splitterG12ton340n421 , splittern251ton421G2570 , 0 , 1 , n421 );
and_AQFP n422_( clk_4 , buf_n420_n422_1 , n421 , 0 , 1 , n422 );
and_AQFP n423_( clk_6 , splitterfromG132 , n422 , 0 , 1 , n423 );
or_AQFP n424_( clk_8 , n419 , n423 , 0 , 0 , n424 );
or_AQFP n425_( clk_1 , n418 , n424 , 0 , 0 , n425 );
or_AQFP n426_( clk_2 , n415 , n425 , 0 , 0 , n426 );
or_AQFP n427_( clk_3 , n385 , n426 , 0 , 0 , n427 );
or_AQFP n428_( clk_5 , n351 , n427 , 0 , 0 , n428 );
and_AQFP n429_( clk_6 , splitterG117ton224n429 , buf_G41_n429_1 , 0 , 1 , n429 );
and_AQFP n430_( clk_5 , splitterG117ton260n429 , buf_G73_n430_1 , 0 , 1 , n430 );
or_AQFP n431_( clk_6 , splitterG120ton240n431 , n430 , 0 , 0 , n431 );
and_AQFP n432_( clk_8 , n429 , n431 , 0 , 1 , n432 );
and_AQFP n433_( clk_7 , buf_G51_n433_1 , splittern203ton272n434 , 0 , 1 , n433 );
and_AQFP n434_( clk_7 , buf_G62_n434_1 , splittern203ton272n434 , 0 , 1 , n434 );
or_AQFP n435_( clk_8 , n433 , n434 , 0 , 0 , n435 );
and_AQFP n436_( clk_2 , n432 , n435 , 0 , 1 , n436 );
and_AQFP n437_( clk_8 , splitterG122ton437n438 , splitterfromn436 , 0 , 1 , n437 );
or_AQFP n438_( clk_2 , splitterG122ton282n438 , n437 , 0 , 0 , n438 );
or_AQFP n439_( clk_4 , splittern191ton330G2558 , splittern294ton408n440 , 0 , 0 , n439 );
and_AQFP n440_( clk_4 , splittern191ton330G2558 , splittern294ton408n440 , 0 , 1 , n440 );
and_AQFP n441_( clk_5 , n439 , n440 , 0 , 1 , n441 );
or_AQFP n442_( clk_7 , splittern184ton442G2557 , splitterfromn441 , 0 , 0 , n442 );
and_AQFP n443_( clk_7 , splittern184ton442G2557 , splitterfromn441 , 1 , 0 , n443 );
and_AQFP n444_( clk_8 , n442 , n443 , 0 , 1 , n444 );
or_AQFP n445_( clk_1 , buf_G29_n445_1 , n444 , 0 , 0 , n445 );
and_AQFP n446_( clk_5 , splitterG123ton446n447 , buf_splitterfromn436_n446_1 , 0 , 1 , n446 );
or_AQFP n447_( clk_6 , splitterG123ton446n447 , n446 , 0 , 0 , n447 );
or_AQFP n448_( clk_1 , buf_G127_n448_1 , splittern198ton325G2559 , 0 , 0 , n448 );
or_AQFP n449_( clk_1 , buf_G30_n449_1 , splittern184ton345G2557 , 0 , 0 , n449 );
or_AQFP n450_( clk_3 , splitterfromn448 , splitterfromn449 , 0 , 0 , n450 );
and_AQFP n451_( clk_6 , splitterG8ton451n486 , splittern450ton451n469 , 1 , 0 , n451 );
and_AQFP n452_( clk_8 , buf_splitterfromG133_n452_1 , splittern451ton452n487 , 1 , 0 , n452 );
or_AQFP n453_( clk_6 , splitterG8ton451n486 , splittern450ton451n469 , 0 , 0 , n453 );
or_AQFP n454_( clk_4 , splittern259ton454G2571 , splittern453ton493n454 , 0 , 0 , n454 );
and_AQFP n455_( clk_8 , buf_splitterfromG132_n455_1 , splittern451ton452n487 , 1 , 0 , n455 );
and_AQFP n456_( clk_7 , buf_splitterfromG129_n456_1 , splittern450ton456n469 , 0 , 0 , n456 );
and_AQFP n457_( clk_7 , buf_splitterG140ton327n457_n457_1 , splittern450ton456n469 , 0 , 1 , n457 );
and_AQFP n458_( clk_8 , n456 , n457 , 0 , 1 , n458 );
and_AQFP n459_( clk_2 , splittern223ton459G2567 , n458 , 0 , 1 , n459 );
and_AQFP n460_( clk_5 , splitterfromG128 , splittern450ton460n469 , 1 , 0 , n460 );
and_AQFP n461_( clk_5 , splitterG139ton396n461 , splittern450ton460n469 , 0 , 1 , n461 );
or_AQFP n462_( clk_6 , n460 , n461 , 0 , 0 , n462 );
and_AQFP n463_( clk_2 , splittern245ton474G2566 , splitterfromn462 , 1 , 0 , n463 );
and_AQFP n464_( clk_5 , splitterfromG126 , splittern450ton460n469 , 1 , 0 , n464 );
and_AQFP n465_( clk_6 , splitterG138ton381n465 , splittern450ton451n469 , 0 , 1 , n465 );
or_AQFP n466_( clk_7 , n464 , n465 , 0 , 0 , n466 );
or_AQFP n467_( clk_1 , splittern275ton467n283 , splitterfromn466 , 0 , 0 , n467 );
and_AQFP n468_( clk_7 , buf_splitterfromG125_n468_1 , splittern450ton456n469 , 1 , 0 , n468 );
and_AQFP n469_( clk_7 , buf_splitterG136ton362n469_n469_1 , splittern450ton456n469 , 0 , 1 , n469 );
or_AQFP n470_( clk_8 , n468 , n469 , 0 , 0 , n470 );
and_AQFP n471_( clk_1 , splittern231ton471n232 , n470 , 1 , 0 , n471 );
and_AQFP n472_( clk_2 , n467 , n471 , 0 , 0 , n472 );
and_AQFP n473_( clk_1 , splittern275ton467n283 , splitterfromn466 , 0 , 0 , n473 );
and_AQFP n474_( clk_1 , splittern245ton474G2566 , splitterfromn462 , 0 , 0 , n474 );
or_AQFP n475_( clk_2 , n473 , n474 , 0 , 0 , n475 );
or_AQFP n476_( clk_3 , n472 , n475 , 0 , 0 , n476 );
and_AQFP n477_( clk_4 , n463 , n476 , 1 , 0 , n477 );
or_AQFP n478_( clk_5 , splitterfromn459 , n477 , 0 , 0 , n478 );
and_AQFP n479_( clk_8 , splitterG8ton479n486 , splittern215ton479G2568 , 0 , 1 , n479 );
and_AQFP n480_( clk_8 , buf_splitterfromG130_n480_1 , splittern451ton452n487 , 0 , 0 , n480 );
and_AQFP n481_( clk_8 , buf_splitterG141ton158n481_n481_1 , splittern453ton481n454 , 0 , 1 , n481 );
and_AQFP n482_( clk_1 , n480 , n481 , 0 , 1 , n482 );
and_AQFP n483_( clk_2 , n479 , n482 , 0 , 1 , n483 );
or_AQFP n484_( clk_4 , splitterfromn459 , splitterfromn483 , 0 , 0 , n484 );
and_AQFP n485_( clk_6 , n478 , n484 , 0 , 1 , n485 );
and_AQFP n486_( clk_8 , splitterG8ton479n486 , splittern207ton486G2569 , 0 , 1 , n486 );
and_AQFP n487_( clk_8 , buf_splitterG131ton368n487_n487_1 , splittern451ton452n487 , 0 , 0 , n487 );
and_AQFP n488_( clk_8 , buf_splitterG142ton332n488_n488_1 , splittern453ton481n454 , 0 , 1 , n488 );
and_AQFP n489_( clk_1 , n487 , n488 , 0 , 1 , n489 );
and_AQFP n490_( clk_2 , n486 , n489 , 0 , 1 , n490 );
or_AQFP n491_( clk_5 , splitterfromn483 , splitterfromn490 , 0 , 0 , n491 );
or_AQFP n492_( clk_7 , n485 , n491 , 0 , 0 , n492 );
and_AQFP n493_( clk_4 , splittern251ton493G2570 , splittern453ton493n454 , 0 , 1 , n493 );
or_AQFP n494_( clk_6 , splitterfromn490 , n493 , 0 , 0 , n494 );
and_AQFP n495_( clk_8 , n492 , n494 , 0 , 1 , n495 );
or_AQFP n496_( clk_1 , buf_n455_n496_1 , n495 , 0 , 0 , n496 );
and_AQFP n497_( clk_2 , buf_n454_n497_1 , n496 , 0 , 0 , n497 );
or_AQFP n498_( clk_3 , buf_n452_n498_1 , n497 , 0 , 0 , n498 );
and_AQFP n499_( clk_3 , splitterfromn448 , splitterfromn449 , 0 , 1 , n499 );
or_AQFP n500_( clk_3 , splitterG136ton500n469 , splitterfromn359 , 0 , 0 , n500 );
and_AQFP n501_( clk_7 , splittern499ton503n512 , splitterfromn500 , 0 , 1 , n501 );
or_AQFP n502_( clk_4 , splitterG138ton502n465 , splitterfromn378 , 0 , 0 , n502 );
and_AQFP n503_( clk_6 , splittern499ton503n512 , n502 , 0 , 1 , n503 );
and_AQFP n504_( clk_1 , n501 , splittern503ton504n522 , 0 , 1 , n504 );
or_AQFP n505_( clk_3 , splitterG135ton505n309 , splittern306ton307n510 , 0 , 0 , n505 );
and_AQFP n506_( clk_4 , splitterG134ton506n401 , splittern267ton399G2572 , 0 , 1 , n506 );
and_AQFP n507_( clk_6 , splitterfromn505 , n506 , 0 , 1 , n507 );
and_AQFP n508_( clk_7 , splittern499ton503n512 , n507 , 0 , 1 , n508 );
or_AQFP n509_( clk_1 , splittern503ton504n522 , n508 , 0 , 0 , n509 );
and_AQFP n510_( clk_4 , splitterG135ton510n309 , splittern306ton307n510 , 0 , 1 , n510 );
and_AQFP n511_( clk_6 , splitterfromn500 , n510 , 0 , 1 , n511 );
and_AQFP n512_( clk_7 , splittern499ton503n512 , n511 , 0 , 1 , n512 );
or_AQFP n513_( clk_3 , splitterG134ton513n401 , splittern267ton399G2572 , 0 , 0 , n513 );
and_AQFP n514_( clk_5 , splittern499ton514n512 , n513 , 0 , 1 , n514 );
or_AQFP n515_( clk_1 , splitterfromn512 , splitterfromn514 , 0 , 0 , n515 );
or_AQFP n516_( clk_3 , n509 , n515 , 0 , 0 , n516 );
and_AQFP n517_( clk_5 , splitterfromn504 , n516 , 0 , 1 , n517 );
and_AQFP n518_( clk_4 , n498 , buf_n517_n518_1 , 0 , 0 , n518 );
and_AQFP n519_( clk_8 , buf_splitterfromn505_n519_1 , splitterfromn514 , 0 , 1 , n519 );
and_AQFP n520_( clk_2 , splitterfromn512 , n519 , 0 , 1 , n520 );
and_AQFP n521_( clk_4 , splitterfromn504 , n520 , 0 , 1 , n521 );
or_AQFP n522_( clk_5 , buf_splittern503ton504n522_n522_1 , n521 , 0 , 0 , n522 );
or_AQFP n523_( clk_5 , n518 , buf_n522_n523_1 , 0 , 0 , n523 );
and_AQFP n524_( clk_3 , splitterfromG10 , splittern176ton524G2556 , 0 , 1 , n524 );
and_AQFP n525_( clk_4 , splitterfromn445 , n524 , 0 , 0 , n525 );
PO_AQFP G2531_( clk_6 , splitterG115toG2531G2549 , 0 , G2531 );
PO_AQFP G2532_( clk_6 , splitterG115toG2531G2549 , 0 , G2532 );
PO_AQFP G2533_( clk_6 , splitterG115toG2531G2549 , 0 , G2533 );
PO_AQFP G2534_( clk_6 , splitterfromG124 , 0 , G2534 );
PO_AQFP G2535_( clk_6 , splitterfromG124 , 0 , G2535 );
PO_AQFP G2536_( clk_6 , splitterG137toG2536G2538 , 0 , G2536 );
PO_AQFP G2537_( clk_6 , splitterG137toG2536G2538 , 0 , G2537 );
PO_AQFP G2538_( clk_6 , splitterG137toG2536G2538 , 0 , G2538 );
PO_AQFP G2539_( clk_6 , buf_splitterfromG32_G2539_1 , 0 , G2539 );
PO_AQFP G2540_( clk_6 , buf_splitterfromG106_G2540_1 , 0 , G2540 );
PO_AQFP G2541_( clk_6 , buf_splitterfromG64_G2541_1 , 0 , G2541 );
PO_AQFP G2542_( clk_6 , buf_splitterfromG76_G2542_1 , 0 , G2542 );
PO_AQFP G2543_( clk_6 , buf_splitterfromG53_G2543_1 , 0 , G2543 );
PO_AQFP G2544_( clk_6 , buf_splitterfromG96_G2544_1 , 0 , G2544 );
PO_AQFP G2545_( clk_6 , buf_splitterfromG43_G2545_1 , 0 , G2545 );
PO_AQFP G2546_( clk_6 , buf_splitterfromG86_G2546_1 , 0 , G2546 );
PO_AQFP G2547_( clk_6 , buf_n160_G2547_1 , 0 , G2547 );
PO_AQFP G2548_( clk_6 , buf_n162_G2548_1 , 0 , G2548 );
PO_AQFP G2549_( clk_6 , splitterG115toG2531G2549 , 0 , G2549 );
PO_AQFP G2550_( clk_6 , buf_n163_G2550_1 , 0 , G2550 );
PO_AQFP G2551_( clk_6 , buf_splittern164ton165G2551_G2551_1 , 0 , G2551 );
PO_AQFP G2552_( clk_6 , buf_n165_G2552_1 , 0 , G2552 );
PO_AQFP G2553_( clk_6 , buf_n166_G2553_1 , 0 , G2553 );
PO_AQFP G2554_( clk_6 , splitterfromn173 , 0 , G2554 );
PO_AQFP G2555_( clk_6 , splitterfromn173 , 0 , G2555 );
PO_AQFP G2556_( clk_6 , buf_splittern176ton524G2556_G2556_1 , 0 , G2556 );
PO_AQFP G2557_( clk_6 , buf_splittern184ton442G2557_G2557_1 , 0 , G2557 );
PO_AQFP G2558_( clk_6 , buf_splittern191ton330G2558_G2558_1 , 0 , G2558 );
PO_AQFP G2559_( clk_6 , buf_splittern198ton325G2559_G2559_1 , 0 , G2559 );
PO_AQFP G2560_( clk_6 , splittern207toG2560G2569 , 0 , G2560 );
PO_AQFP G2561_( clk_6 , splittern215toG2561G2568 , 0 , G2561 );
PO_AQFP G2562_( clk_6 , splittern223toG2562G2567 , 0 , G2562 );
PO_AQFP G2563_( clk_6 , buf_n232_G2563_1 , 0 , G2563 );
PO_AQFP G2564_( clk_6 , n235 , 0 , G2564 );
PO_AQFP G2565_( clk_6 , buf_n237_G2565_1 , 0 , G2565 );
PO_AQFP G2566_( clk_6 , buf_splittern245ton279G2566_G2566_1 , 0 , G2566 );
PO_AQFP G2567_( clk_6 , splittern223toG2562G2567 , 0 , G2567 );
PO_AQFP G2568_( clk_6 , splittern215toG2561G2568 , 0 , G2568 );
PO_AQFP G2569_( clk_6 , splittern207toG2560G2569 , 0 , G2569 );
PO_AQFP G2570_( clk_6 , buf_splittern251ton493G2570_G2570_1 , 0 , G2570 );
PO_AQFP G2571_( clk_6 , buf_splittern259ton454G2571_G2571_1 , 0 , G2571 );
PO_AQFP G2572_( clk_6 , buf_splittern267ton399G2572_G2572_1 , 0 , G2572 );
PO_AQFP G2573_( clk_6 , splitterfromn278 , 0 , G2573 );
PO_AQFP G2574_( clk_6 , splitterfromn278 , 0 , G2574 );
PO_AQFP G2575_( clk_6 , splitterfromn281 , 0 , G2575 );
PO_AQFP G2576_( clk_6 , splitterfromn281 , 0 , G2576 );
PO_AQFP G2577_( clk_6 , buf_n283_G2577_1 , 0 , G2577 );
PO_AQFP G2578_( clk_6 , splitterfromn287 , 0 , G2578 );
PO_AQFP G2579_( clk_6 , splitterfromn287 , 0 , G2579 );
PO_AQFP G2580_( clk_6 , buf_n298_G2580_1 , 0 , G2580 );
PO_AQFP G2581_( clk_6 , buf_splitterfromG10_G2581_1 , 1 , G2581 );
PO_AQFP G2584_( clk_6 , splitterfromn428 , 0 , G2584 );
PO_AQFP G2585_( clk_6 , splitterfromn428 , 0 , G2585 );
PO_AQFP G2586_( clk_6 , buf_n438_G2586_1 , 0 , G2586 );
PO_AQFP G2587_( clk_6 , buf_splitterfromn445_G2587_1 , 0 , G2587 );
PO_AQFP G2588_( clk_6 , splitterfromn447 , 0 , G2588 );
PO_AQFP G2589_( clk_6 , splitterfromn447 , 0 , G2589 );
PO_AQFP G2591_( clk_6 , n523 , 1 , G2591 );
PO_AQFP G2593_( clk_6 , splitterfromn525 , 1 , G2593 );
PO_AQFP G2594_( clk_6 , splitterfromn525 , 1 , G2594 );
buf_AQFP buf_G10_splitterfromG10_11_( clk_3 , G10 , 0 , buf_G10_splitterfromG10_11 );
buf_AQFP buf_G10_splitterfromG10_10_( clk_5 , buf_G10_splitterfromG10_11 , 0 , buf_G10_splitterfromG10_10 );
buf_AQFP buf_G10_splitterfromG10_9_( clk_7 , buf_G10_splitterfromG10_10 , 0 , buf_G10_splitterfromG10_9 );
buf_AQFP buf_G10_splitterfromG10_8_( clk_1 , buf_G10_splitterfromG10_9 , 0 , buf_G10_splitterfromG10_8 );
buf_AQFP buf_G10_splitterfromG10_7_( clk_3 , buf_G10_splitterfromG10_8 , 0 , buf_G10_splitterfromG10_7 );
buf_AQFP buf_G10_splitterfromG10_6_( clk_5 , buf_G10_splitterfromG10_7 , 0 , buf_G10_splitterfromG10_6 );
buf_AQFP buf_G10_splitterfromG10_5_( clk_7 , buf_G10_splitterfromG10_6 , 0 , buf_G10_splitterfromG10_5 );
buf_AQFP buf_G10_splitterfromG10_4_( clk_1 , buf_G10_splitterfromG10_5 , 0 , buf_G10_splitterfromG10_4 );
buf_AQFP buf_G10_splitterfromG10_3_( clk_3 , buf_G10_splitterfromG10_4 , 0 , buf_G10_splitterfromG10_3 );
buf_AQFP buf_G10_splitterfromG10_2_( clk_5 , buf_G10_splitterfromG10_3 , 0 , buf_G10_splitterfromG10_2 );
buf_AQFP buf_G10_splitterfromG10_1_( clk_7 , buf_G10_splitterfromG10_2 , 0 , buf_G10_splitterfromG10_1 );
buf_AQFP buf_G100_n195_1_( clk_3 , G100 , 0 , buf_G100_n195_1 );
buf_AQFP buf_G101_n388_2_( clk_3 , G101 , 0 , buf_G101_n388_2 );
buf_AQFP buf_G101_n388_1_( clk_5 , buf_G101_n388_2 , 0 , buf_G101_n388_1 );
buf_AQFP buf_G102_n373_2_( clk_3 , G102 , 0 , buf_G102_n373_2 );
buf_AQFP buf_G102_n373_1_( clk_5 , buf_G102_n373_2 , 0 , buf_G102_n373_1 );
buf_AQFP buf_G103_n354_2_( clk_3 , G103 , 0 , buf_G103_n354_2 );
buf_AQFP buf_G103_n354_1_( clk_5 , buf_G103_n354_2 , 0 , buf_G103_n354_1 );
buf_AQFP buf_G105_n304_2_( clk_3 , G105 , 0 , buf_G105_n304_2 );
buf_AQFP buf_G105_n304_1_( clk_5 , buf_G105_n304_2 , 0 , buf_G105_n304_1 );
buf_AQFP buf_G106_splitterfromG106_7_( clk_3 , G106 , 0 , buf_G106_splitterfromG106_7 );
buf_AQFP buf_G106_splitterfromG106_6_( clk_5 , buf_G106_splitterfromG106_7 , 0 , buf_G106_splitterfromG106_6 );
buf_AQFP buf_G106_splitterfromG106_5_( clk_7 , buf_G106_splitterfromG106_6 , 0 , buf_G106_splitterfromG106_5 );
buf_AQFP buf_G106_splitterfromG106_4_( clk_1 , buf_G106_splitterfromG106_5 , 0 , buf_G106_splitterfromG106_4 );
buf_AQFP buf_G106_splitterfromG106_3_( clk_3 , buf_G106_splitterfromG106_4 , 0 , buf_G106_splitterfromG106_3 );
buf_AQFP buf_G106_splitterfromG106_2_( clk_5 , buf_G106_splitterfromG106_3 , 0 , buf_G106_splitterfromG106_2 );
buf_AQFP buf_G106_splitterfromG106_1_( clk_7 , buf_G106_splitterfromG106_2 , 0 , buf_G106_splitterfromG106_1 );
buf_AQFP buf_G107_n291_2_( clk_3 , G107 , 0 , buf_G107_n291_2 );
buf_AQFP buf_G107_n291_1_( clk_5 , buf_G107_n291_2 , 0 , buf_G107_n291_1 );
buf_AQFP buf_G108_n185_2_( clk_3 , G108 , 0 , buf_G108_n185_2 );
buf_AQFP buf_G108_n185_1_( clk_5 , buf_G108_n185_2 , 0 , buf_G108_n185_1 );
buf_AQFP buf_G109_n178_1_( clk_3 , G109 , 0 , buf_G109_n178_1 );
buf_AQFP buf_G11_n162_1_( clk_3 , G11 , 0 , buf_G11_n162_1 );
buf_AQFP buf_G110_n196_1_( clk_3 , G110 , 0 , buf_G110_n196_1 );
buf_AQFP buf_G111_n390_2_( clk_3 , G111 , 0 , buf_G111_n390_2 );
buf_AQFP buf_G111_n390_1_( clk_5 , buf_G111_n390_2 , 0 , buf_G111_n390_1 );
buf_AQFP buf_G112_n375_2_( clk_3 , G112 , 0 , buf_G112_n375_2 );
buf_AQFP buf_G112_n375_1_( clk_5 , buf_G112_n375_2 , 0 , buf_G112_n375_1 );
buf_AQFP buf_G113_n356_2_( clk_3 , G113 , 0 , buf_G113_n356_2 );
buf_AQFP buf_G113_n356_1_( clk_5 , buf_G113_n356_2 , 0 , buf_G113_n356_1 );
buf_AQFP buf_G116_n233_1_( clk_3 , G116 , 0 , buf_G116_n233_1 );
buf_AQFP buf_G118_splitterfromG118_5_( clk_3 , G118 , 0 , buf_G118_splitterfromG118_5 );
buf_AQFP buf_G118_splitterfromG118_4_( clk_5 , buf_G118_splitterfromG118_5 , 0 , buf_G118_splitterfromG118_4 );
buf_AQFP buf_G118_splitterfromG118_3_( clk_7 , buf_G118_splitterfromG118_4 , 0 , buf_G118_splitterfromG118_3 );
buf_AQFP buf_G118_splitterfromG118_2_( clk_1 , buf_G118_splitterfromG118_3 , 0 , buf_G118_splitterfromG118_2 );
buf_AQFP buf_G118_splitterfromG118_1_( clk_3 , buf_G118_splitterfromG118_2 , 0 , buf_G118_splitterfromG118_1 );
buf_AQFP buf_G119_splitterfromG119_9_( clk_3 , G119 , 0 , buf_G119_splitterfromG119_9 );
buf_AQFP buf_G119_splitterfromG119_8_( clk_5 , buf_G119_splitterfromG119_9 , 0 , buf_G119_splitterfromG119_8 );
buf_AQFP buf_G119_splitterfromG119_7_( clk_7 , buf_G119_splitterfromG119_8 , 0 , buf_G119_splitterfromG119_7 );
buf_AQFP buf_G119_splitterfromG119_6_( clk_1 , buf_G119_splitterfromG119_7 , 0 , buf_G119_splitterfromG119_6 );
buf_AQFP buf_G119_splitterfromG119_5_( clk_3 , buf_G119_splitterfromG119_6 , 0 , buf_G119_splitterfromG119_5 );
buf_AQFP buf_G119_splitterfromG119_4_( clk_5 , buf_G119_splitterfromG119_5 , 0 , buf_G119_splitterfromG119_4 );
buf_AQFP buf_G119_splitterfromG119_3_( clk_7 , buf_G119_splitterfromG119_4 , 0 , buf_G119_splitterfromG119_3 );
buf_AQFP buf_G119_splitterfromG119_2_( clk_1 , buf_G119_splitterfromG119_3 , 0 , buf_G119_splitterfromG119_2 );
buf_AQFP buf_G119_splitterfromG119_1_( clk_3 , buf_G119_splitterfromG119_2 , 0 , buf_G119_splitterfromG119_1 );
buf_AQFP buf_G122_splitterG122ton437n438_6_( clk_3 , G122 , 0 , buf_G122_splitterG122ton437n438_6 );
buf_AQFP buf_G122_splitterG122ton437n438_5_( clk_5 , buf_G122_splitterG122ton437n438_6 , 0 , buf_G122_splitterG122ton437n438_5 );
buf_AQFP buf_G122_splitterG122ton437n438_4_( clk_7 , buf_G122_splitterG122ton437n438_5 , 0 , buf_G122_splitterG122ton437n438_4 );
buf_AQFP buf_G122_splitterG122ton437n438_3_( clk_1 , buf_G122_splitterG122ton437n438_4 , 0 , buf_G122_splitterG122ton437n438_3 );
buf_AQFP buf_G122_splitterG122ton437n438_2_( clk_3 , buf_G122_splitterG122ton437n438_3 , 0 , buf_G122_splitterG122ton437n438_2 );
buf_AQFP buf_G122_splitterG122ton437n438_1_( clk_5 , buf_G122_splitterG122ton437n438_2 , 0 , buf_G122_splitterG122ton437n438_1 );
buf_AQFP buf_G123_splitterG123ton285n447_5_( clk_3 , G123 , 0 , buf_G123_splitterG123ton285n447_5 );
buf_AQFP buf_G123_splitterG123ton285n447_4_( clk_5 , buf_G123_splitterG123ton285n447_5 , 0 , buf_G123_splitterG123ton285n447_4 );
buf_AQFP buf_G123_splitterG123ton285n447_3_( clk_7 , buf_G123_splitterG123ton285n447_4 , 0 , buf_G123_splitterG123ton285n447_3 );
buf_AQFP buf_G123_splitterG123ton285n447_2_( clk_1 , buf_G123_splitterG123ton285n447_3 , 0 , buf_G123_splitterG123ton285n447_2 );
buf_AQFP buf_G123_splitterG123ton285n447_1_( clk_3 , buf_G123_splitterG123ton285n447_2 , 0 , buf_G123_splitterG123ton285n447_1 );
buf_AQFP buf_G124_splitterfromG124_13_( clk_3 , G124 , 0 , buf_G124_splitterfromG124_13 );
buf_AQFP buf_G124_splitterfromG124_12_( clk_5 , buf_G124_splitterfromG124_13 , 0 , buf_G124_splitterfromG124_12 );
buf_AQFP buf_G124_splitterfromG124_11_( clk_7 , buf_G124_splitterfromG124_12 , 0 , buf_G124_splitterfromG124_11 );
buf_AQFP buf_G124_splitterfromG124_10_( clk_1 , buf_G124_splitterfromG124_11 , 0 , buf_G124_splitterfromG124_10 );
buf_AQFP buf_G124_splitterfromG124_9_( clk_3 , buf_G124_splitterfromG124_10 , 0 , buf_G124_splitterfromG124_9 );
buf_AQFP buf_G124_splitterfromG124_8_( clk_5 , buf_G124_splitterfromG124_9 , 0 , buf_G124_splitterfromG124_8 );
buf_AQFP buf_G124_splitterfromG124_7_( clk_7 , buf_G124_splitterfromG124_8 , 0 , buf_G124_splitterfromG124_7 );
buf_AQFP buf_G124_splitterfromG124_6_( clk_1 , buf_G124_splitterfromG124_7 , 0 , buf_G124_splitterfromG124_6 );
buf_AQFP buf_G124_splitterfromG124_5_( clk_3 , buf_G124_splitterfromG124_6 , 0 , buf_G124_splitterfromG124_5 );
buf_AQFP buf_G124_splitterfromG124_4_( clk_5 , buf_G124_splitterfromG124_5 , 0 , buf_G124_splitterfromG124_4 );
buf_AQFP buf_G124_splitterfromG124_3_( clk_7 , buf_G124_splitterfromG124_4 , 0 , buf_G124_splitterfromG124_3 );
buf_AQFP buf_G124_splitterfromG124_2_( clk_1 , buf_G124_splitterfromG124_3 , 0 , buf_G124_splitterfromG124_2 );
buf_AQFP buf_G124_splitterfromG124_1_( clk_3 , buf_G124_splitterfromG124_2 , 0 , buf_G124_splitterfromG124_1 );
buf_AQFP buf_G125_splitterfromG125_5_( clk_3 , G125 , 0 , buf_G125_splitterfromG125_5 );
buf_AQFP buf_G125_splitterfromG125_4_( clk_5 , buf_G125_splitterfromG125_5 , 0 , buf_G125_splitterfromG125_4 );
buf_AQFP buf_G125_splitterfromG125_3_( clk_7 , buf_G125_splitterfromG125_4 , 0 , buf_G125_splitterfromG125_3 );
buf_AQFP buf_G125_splitterfromG125_2_( clk_1 , buf_G125_splitterfromG125_3 , 0 , buf_G125_splitterfromG125_2 );
buf_AQFP buf_G125_splitterfromG125_1_( clk_3 , buf_G125_splitterfromG125_2 , 0 , buf_G125_splitterfromG125_1 );
buf_AQFP buf_G126_splitterfromG126_4_( clk_3 , G126 , 0 , buf_G126_splitterfromG126_4 );
buf_AQFP buf_G126_splitterfromG126_3_( clk_5 , buf_G126_splitterfromG126_4 , 0 , buf_G126_splitterfromG126_3 );
buf_AQFP buf_G126_splitterfromG126_2_( clk_7 , buf_G126_splitterfromG126_3 , 0 , buf_G126_splitterfromG126_2 );
buf_AQFP buf_G126_splitterfromG126_1_( clk_1 , buf_G126_splitterfromG126_2 , 0 , buf_G126_splitterfromG126_1 );
buf_AQFP buf_G127_n448_3_( clk_3 , G127 , 0 , buf_G127_n448_3 );
buf_AQFP buf_G127_n448_2_( clk_5 , buf_G127_n448_3 , 0 , buf_G127_n448_2 );
buf_AQFP buf_G127_n448_1_( clk_7 , buf_G127_n448_2 , 0 , buf_G127_n448_1 );
buf_AQFP buf_G128_splitterfromG128_4_( clk_3 , G128 , 0 , buf_G128_splitterfromG128_4 );
buf_AQFP buf_G128_splitterfromG128_3_( clk_5 , buf_G128_splitterfromG128_4 , 0 , buf_G128_splitterfromG128_3 );
buf_AQFP buf_G128_splitterfromG128_2_( clk_7 , buf_G128_splitterfromG128_3 , 0 , buf_G128_splitterfromG128_2 );
buf_AQFP buf_G128_splitterfromG128_1_( clk_1 , buf_G128_splitterfromG128_2 , 0 , buf_G128_splitterfromG128_1 );
buf_AQFP buf_G129_splitterfromG129_4_( clk_3 , G129 , 0 , buf_G129_splitterfromG129_4 );
buf_AQFP buf_G129_splitterfromG129_3_( clk_5 , buf_G129_splitterfromG129_4 , 0 , buf_G129_splitterfromG129_3 );
buf_AQFP buf_G129_splitterfromG129_2_( clk_7 , buf_G129_splitterfromG129_3 , 0 , buf_G129_splitterfromG129_2 );
buf_AQFP buf_G129_splitterfromG129_1_( clk_1 , buf_G129_splitterfromG129_2 , 0 , buf_G129_splitterfromG129_1 );
buf_AQFP buf_G130_splitterfromG130_4_( clk_3 , G130 , 0 , buf_G130_splitterfromG130_4 );
buf_AQFP buf_G130_splitterfromG130_3_( clk_5 , buf_G130_splitterfromG130_4 , 0 , buf_G130_splitterfromG130_3 );
buf_AQFP buf_G130_splitterfromG130_2_( clk_7 , buf_G130_splitterfromG130_3 , 0 , buf_G130_splitterfromG130_2 );
buf_AQFP buf_G130_splitterfromG130_1_( clk_1 , buf_G130_splitterfromG130_2 , 0 , buf_G130_splitterfromG130_1 );
buf_AQFP buf_G131_splitterG131ton368n487_5_( clk_3 , G131 , 0 , buf_G131_splitterG131ton368n487_5 );
buf_AQFP buf_G131_splitterG131ton368n487_4_( clk_5 , buf_G131_splitterG131ton368n487_5 , 0 , buf_G131_splitterG131ton368n487_4 );
buf_AQFP buf_G131_splitterG131ton368n487_3_( clk_7 , buf_G131_splitterG131ton368n487_4 , 0 , buf_G131_splitterG131ton368n487_3 );
buf_AQFP buf_G131_splitterG131ton368n487_2_( clk_1 , buf_G131_splitterG131ton368n487_3 , 0 , buf_G131_splitterG131ton368n487_2 );
buf_AQFP buf_G131_splitterG131ton368n487_1_( clk_3 , buf_G131_splitterG131ton368n487_2 , 0 , buf_G131_splitterG131ton368n487_1 );
buf_AQFP buf_G132_splitterfromG132_5_( clk_3 , G132 , 0 , buf_G132_splitterfromG132_5 );
buf_AQFP buf_G132_splitterfromG132_4_( clk_5 , buf_G132_splitterfromG132_5 , 0 , buf_G132_splitterfromG132_4 );
buf_AQFP buf_G132_splitterfromG132_3_( clk_7 , buf_G132_splitterfromG132_4 , 0 , buf_G132_splitterfromG132_3 );
buf_AQFP buf_G132_splitterfromG132_2_( clk_1 , buf_G132_splitterfromG132_3 , 0 , buf_G132_splitterfromG132_2 );
buf_AQFP buf_G132_splitterfromG132_1_( clk_3 , buf_G132_splitterfromG132_2 , 0 , buf_G132_splitterfromG132_1 );
buf_AQFP buf_G133_splitterfromG133_5_( clk_3 , G133 , 0 , buf_G133_splitterfromG133_5 );
buf_AQFP buf_G133_splitterfromG133_4_( clk_5 , buf_G133_splitterfromG133_5 , 0 , buf_G133_splitterfromG133_4 );
buf_AQFP buf_G133_splitterfromG133_3_( clk_7 , buf_G133_splitterfromG133_4 , 0 , buf_G133_splitterfromG133_3 );
buf_AQFP buf_G133_splitterfromG133_2_( clk_1 , buf_G133_splitterfromG133_3 , 0 , buf_G133_splitterfromG133_2 );
buf_AQFP buf_G133_splitterfromG133_1_( clk_3 , buf_G133_splitterfromG133_2 , 0 , buf_G133_splitterfromG133_1 );
buf_AQFP buf_G134_splitterG134ton513n401_3_( clk_3 , G134 , 0 , buf_G134_splitterG134ton513n401_3 );
buf_AQFP buf_G134_splitterG134ton513n401_2_( clk_5 , buf_G134_splitterG134ton513n401_3 , 0 , buf_G134_splitterG134ton513n401_2 );
buf_AQFP buf_G134_splitterG134ton513n401_1_( clk_7 , buf_G134_splitterG134ton513n401_2 , 0 , buf_G134_splitterG134ton513n401_1 );
buf_AQFP buf_G135_splitterG135ton505n309_3_( clk_3 , G135 , 0 , buf_G135_splitterG135ton505n309_3 );
buf_AQFP buf_G135_splitterG135ton505n309_2_( clk_5 , buf_G135_splitterG135ton505n309_3 , 0 , buf_G135_splitterG135ton505n309_2 );
buf_AQFP buf_G135_splitterG135ton505n309_1_( clk_7 , buf_G135_splitterG135ton505n309_2 , 0 , buf_G135_splitterG135ton505n309_1 );
buf_AQFP buf_G136_splitterG136ton500n469_3_( clk_3 , G136 , 0 , buf_G136_splitterG136ton500n469_3 );
buf_AQFP buf_G136_splitterG136ton500n469_2_( clk_5 , buf_G136_splitterG136ton500n469_3 , 0 , buf_G136_splitterG136ton500n469_2 );
buf_AQFP buf_G136_splitterG136ton500n469_1_( clk_7 , buf_G136_splitterG136ton500n469_2 , 0 , buf_G136_splitterG136ton500n469_1 );
buf_AQFP buf_G137_splitterG137toG2536G2538_13_( clk_3 , G137 , 0 , buf_G137_splitterG137toG2536G2538_13 );
buf_AQFP buf_G137_splitterG137toG2536G2538_12_( clk_5 , buf_G137_splitterG137toG2536G2538_13 , 0 , buf_G137_splitterG137toG2536G2538_12 );
buf_AQFP buf_G137_splitterG137toG2536G2538_11_( clk_7 , buf_G137_splitterG137toG2536G2538_12 , 0 , buf_G137_splitterG137toG2536G2538_11 );
buf_AQFP buf_G137_splitterG137toG2536G2538_10_( clk_1 , buf_G137_splitterG137toG2536G2538_11 , 0 , buf_G137_splitterG137toG2536G2538_10 );
buf_AQFP buf_G137_splitterG137toG2536G2538_9_( clk_3 , buf_G137_splitterG137toG2536G2538_10 , 0 , buf_G137_splitterG137toG2536G2538_9 );
buf_AQFP buf_G137_splitterG137toG2536G2538_8_( clk_5 , buf_G137_splitterG137toG2536G2538_9 , 0 , buf_G137_splitterG137toG2536G2538_8 );
buf_AQFP buf_G137_splitterG137toG2536G2538_7_( clk_7 , buf_G137_splitterG137toG2536G2538_8 , 0 , buf_G137_splitterG137toG2536G2538_7 );
buf_AQFP buf_G137_splitterG137toG2536G2538_6_( clk_1 , buf_G137_splitterG137toG2536G2538_7 , 0 , buf_G137_splitterG137toG2536G2538_6 );
buf_AQFP buf_G137_splitterG137toG2536G2538_5_( clk_3 , buf_G137_splitterG137toG2536G2538_6 , 0 , buf_G137_splitterG137toG2536G2538_5 );
buf_AQFP buf_G137_splitterG137toG2536G2538_4_( clk_5 , buf_G137_splitterG137toG2536G2538_5 , 0 , buf_G137_splitterG137toG2536G2538_4 );
buf_AQFP buf_G137_splitterG137toG2536G2538_3_( clk_7 , buf_G137_splitterG137toG2536G2538_4 , 0 , buf_G137_splitterG137toG2536G2538_3 );
buf_AQFP buf_G137_splitterG137toG2536G2538_2_( clk_1 , buf_G137_splitterG137toG2536G2538_3 , 0 , buf_G137_splitterG137toG2536G2538_2 );
buf_AQFP buf_G137_splitterG137toG2536G2538_1_( clk_3 , buf_G137_splitterG137toG2536G2538_2 , 0 , buf_G137_splitterG137toG2536G2538_1 );
buf_AQFP buf_G138_splitterG138ton502n465_4_( clk_3 , G138 , 0 , buf_G138_splitterG138ton502n465_4 );
buf_AQFP buf_G138_splitterG138ton502n465_3_( clk_5 , buf_G138_splitterG138ton502n465_4 , 0 , buf_G138_splitterG138ton502n465_3 );
buf_AQFP buf_G138_splitterG138ton502n465_2_( clk_7 , buf_G138_splitterG138ton502n465_3 , 0 , buf_G138_splitterG138ton502n465_2 );
buf_AQFP buf_G138_splitterG138ton502n465_1_( clk_1 , buf_G138_splitterG138ton502n465_2 , 0 , buf_G138_splitterG138ton502n465_1 );
buf_AQFP buf_G139_splitterG139ton159n461_3_( clk_3 , G139 , 0 , buf_G139_splitterG139ton159n461_3 );
buf_AQFP buf_G139_splitterG139ton159n461_2_( clk_5 , buf_G139_splitterG139ton159n461_3 , 0 , buf_G139_splitterG139ton159n461_2 );
buf_AQFP buf_G139_splitterG139ton159n461_1_( clk_7 , buf_G139_splitterG139ton159n461_2 , 0 , buf_G139_splitterG139ton159n461_1 );
buf_AQFP buf_G14_n335_2_( clk_3 , G14 , 0 , buf_G14_n335_2 );
buf_AQFP buf_G14_n335_1_( clk_5 , buf_G14_n335_2 , 0 , buf_G14_n335_1 );
buf_AQFP buf_G140_splitterG140ton159n457_3_( clk_3 , G140 , 0 , buf_G140_splitterG140ton159n457_3 );
buf_AQFP buf_G140_splitterG140ton159n457_2_( clk_5 , buf_G140_splitterG140ton159n457_3 , 0 , buf_G140_splitterG140ton159n457_2 );
buf_AQFP buf_G140_splitterG140ton159n457_1_( clk_7 , buf_G140_splitterG140ton159n457_2 , 0 , buf_G140_splitterG140ton159n457_1 );
buf_AQFP buf_G141_splitterG141ton158n481_4_( clk_3 , G141 , 0 , buf_G141_splitterG141ton158n481_4 );
buf_AQFP buf_G141_splitterG141ton158n481_3_( clk_5 , buf_G141_splitterG141ton158n481_4 , 0 , buf_G141_splitterG141ton158n481_3 );
buf_AQFP buf_G141_splitterG141ton158n481_2_( clk_7 , buf_G141_splitterG141ton158n481_3 , 0 , buf_G141_splitterG141ton158n481_2 );
buf_AQFP buf_G141_splitterG141ton158n481_1_( clk_1 , buf_G141_splitterG141ton158n481_2 , 0 , buf_G141_splitterG141ton158n481_1 );
buf_AQFP buf_G142_splitterG142ton158n488_3_( clk_3 , G142 , 0 , buf_G142_splitterG142ton158n488_3 );
buf_AQFP buf_G142_splitterG142ton158n488_2_( clk_5 , buf_G142_splitterG142ton158n488_3 , 0 , buf_G142_splitterG142ton158n488_2 );
buf_AQFP buf_G142_splitterG142ton158n488_1_( clk_7 , buf_G142_splitterG142ton158n488_2 , 0 , buf_G142_splitterG142ton158n488_1 );
buf_AQFP buf_G143_splitterfromG143_3_( clk_3 , G143 , 0 , buf_G143_splitterfromG143_3 );
buf_AQFP buf_G143_splitterfromG143_2_( clk_5 , buf_G143_splitterfromG143_3 , 0 , buf_G143_splitterfromG143_2 );
buf_AQFP buf_G143_splitterfromG143_1_( clk_7 , buf_G143_splitterfromG143_2 , 0 , buf_G143_splitterfromG143_1 );
buf_AQFP buf_G144_n298_5_( clk_3 , G144 , 0 , buf_G144_n298_5 );
buf_AQFP buf_G144_n298_4_( clk_5 , buf_G144_n298_5 , 0 , buf_G144_n298_4 );
buf_AQFP buf_G144_n298_3_( clk_7 , buf_G144_n298_4 , 0 , buf_G144_n298_3 );
buf_AQFP buf_G144_n298_2_( clk_1 , buf_G144_n298_3 , 0 , buf_G144_n298_2 );
buf_AQFP buf_G144_n298_1_( clk_3 , buf_G144_n298_2 , 0 , buf_G144_n298_1 );
buf_AQFP buf_G147_splitterfromG147_9_( clk_3 , G147 , 0 , buf_G147_splitterfromG147_9 );
buf_AQFP buf_G147_splitterfromG147_8_( clk_5 , buf_G147_splitterfromG147_9 , 0 , buf_G147_splitterfromG147_8 );
buf_AQFP buf_G147_splitterfromG147_7_( clk_7 , buf_G147_splitterfromG147_8 , 0 , buf_G147_splitterfromG147_7 );
buf_AQFP buf_G147_splitterfromG147_6_( clk_1 , buf_G147_splitterfromG147_7 , 0 , buf_G147_splitterfromG147_6 );
buf_AQFP buf_G147_splitterfromG147_5_( clk_3 , buf_G147_splitterfromG147_6 , 0 , buf_G147_splitterfromG147_5 );
buf_AQFP buf_G147_splitterfromG147_4_( clk_5 , buf_G147_splitterfromG147_5 , 0 , buf_G147_splitterfromG147_4 );
buf_AQFP buf_G147_splitterfromG147_3_( clk_7 , buf_G147_splitterfromG147_4 , 0 , buf_G147_splitterfromG147_3 );
buf_AQFP buf_G147_splitterfromG147_2_( clk_1 , buf_G147_splitterfromG147_3 , 0 , buf_G147_splitterfromG147_2 );
buf_AQFP buf_G147_splitterfromG147_1_( clk_3 , buf_G147_splitterfromG147_2 , 0 , buf_G147_splitterfromG147_1 );
buf_AQFP buf_G15_n314_1_( clk_3 , G15 , 0 , buf_G15_n314_1 );
buf_AQFP buf_G16_n365_3_( clk_3 , G16 , 0 , buf_G16_n365_3 );
buf_AQFP buf_G16_n365_2_( clk_5 , buf_G16_n365_3 , 0 , buf_G16_n365_2 );
buf_AQFP buf_G16_n365_1_( clk_7 , buf_G16_n365_2 , 0 , buf_G16_n365_1 );
buf_AQFP buf_G17_n420_2_( clk_3 , G17 , 0 , buf_G17_n420_2 );
buf_AQFP buf_G17_n420_1_( clk_5 , buf_G17_n420_2 , 0 , buf_G17_n420_1 );
buf_AQFP buf_G18_n398_2_( clk_3 , G18 , 0 , buf_G18_n398_2 );
buf_AQFP buf_G18_n398_1_( clk_5 , buf_G18_n398_2 , 0 , buf_G18_n398_1 );
buf_AQFP buf_G19_n299_2_( clk_3 , G19 , 0 , buf_G19_n299_2 );
buf_AQFP buf_G19_n299_1_( clk_5 , buf_G19_n299_2 , 0 , buf_G19_n299_1 );
buf_AQFP buf_G20_n371_4_( clk_3 , G20 , 0 , buf_G20_n371_4 );
buf_AQFP buf_G20_n371_3_( clk_5 , buf_G20_n371_4 , 0 , buf_G20_n371_3 );
buf_AQFP buf_G20_n371_2_( clk_7 , buf_G20_n371_3 , 0 , buf_G20_n371_2 );
buf_AQFP buf_G20_n371_1_( clk_1 , buf_G20_n371_2 , 0 , buf_G20_n371_1 );
buf_AQFP buf_G21_n324_2_( clk_3 , G21 , 0 , buf_G21_n324_2 );
buf_AQFP buf_G21_n324_1_( clk_5 , buf_G21_n324_2 , 0 , buf_G21_n324_1 );
buf_AQFP buf_G24_n352_1_( clk_3 , G24 , 0 , buf_G24_n352_1 );
buf_AQFP buf_G25_n386_1_( clk_3 , G25 , 0 , buf_G25_n386_1 );
buf_AQFP buf_G26_n344_3_( clk_3 , G26 , 0 , buf_G26_n344_3 );
buf_AQFP buf_G26_n344_2_( clk_5 , buf_G26_n344_3 , 0 , buf_G26_n344_2 );
buf_AQFP buf_G26_n344_1_( clk_7 , buf_G26_n344_2 , 0 , buf_G26_n344_1 );
buf_AQFP buf_G27_n329_2_( clk_3 , G27 , 0 , buf_G27_n329_2 );
buf_AQFP buf_G27_n329_1_( clk_5 , buf_G27_n329_2 , 0 , buf_G27_n329_1 );
buf_AQFP buf_G28_n235_13_( clk_3 , G28 , 0 , buf_G28_n235_13 );
buf_AQFP buf_G28_n235_12_( clk_5 , buf_G28_n235_13 , 0 , buf_G28_n235_12 );
buf_AQFP buf_G28_n235_11_( clk_7 , buf_G28_n235_12 , 0 , buf_G28_n235_11 );
buf_AQFP buf_G28_n235_10_( clk_1 , buf_G28_n235_11 , 0 , buf_G28_n235_10 );
buf_AQFP buf_G28_n235_9_( clk_3 , buf_G28_n235_10 , 0 , buf_G28_n235_9 );
buf_AQFP buf_G28_n235_8_( clk_5 , buf_G28_n235_9 , 0 , buf_G28_n235_8 );
buf_AQFP buf_G28_n235_7_( clk_7 , buf_G28_n235_8 , 0 , buf_G28_n235_7 );
buf_AQFP buf_G28_n235_6_( clk_1 , buf_G28_n235_7 , 0 , buf_G28_n235_6 );
buf_AQFP buf_G28_n235_5_( clk_3 , buf_G28_n235_6 , 0 , buf_G28_n235_5 );
buf_AQFP buf_G28_n235_4_( clk_5 , buf_G28_n235_5 , 0 , buf_G28_n235_4 );
buf_AQFP buf_G28_n235_3_( clk_7 , buf_G28_n235_4 , 0 , buf_G28_n235_3 );
buf_AQFP buf_G28_n235_2_( clk_1 , buf_G28_n235_3 , 0 , buf_G28_n235_2 );
buf_AQFP buf_G28_n235_1_( clk_3 , buf_G28_n235_2 , 0 , buf_G28_n235_1 );
buf_AQFP buf_G29_n445_7_( clk_3 , G29 , 0 , buf_G29_n445_7 );
buf_AQFP buf_G29_n445_6_( clk_5 , buf_G29_n445_7 , 0 , buf_G29_n445_6 );
buf_AQFP buf_G29_n445_5_( clk_7 , buf_G29_n445_6 , 0 , buf_G29_n445_5 );
buf_AQFP buf_G29_n445_4_( clk_1 , buf_G29_n445_5 , 0 , buf_G29_n445_4 );
buf_AQFP buf_G29_n445_3_( clk_3 , buf_G29_n445_4 , 0 , buf_G29_n445_3 );
buf_AQFP buf_G29_n445_2_( clk_5 , buf_G29_n445_3 , 0 , buf_G29_n445_2 );
buf_AQFP buf_G29_n445_1_( clk_7 , buf_G29_n445_2 , 0 , buf_G29_n445_1 );
buf_AQFP buf_G30_n449_3_( clk_3 , G30 , 0 , buf_G30_n449_3 );
buf_AQFP buf_G30_n449_2_( clk_5 , buf_G30_n449_3 , 0 , buf_G30_n449_2 );
buf_AQFP buf_G30_n449_1_( clk_7 , buf_G30_n449_2 , 0 , buf_G30_n449_1 );
buf_AQFP buf_G31_n224_2_( clk_3 , G31 , 0 , buf_G31_n224_2 );
buf_AQFP buf_G31_n224_1_( clk_5 , buf_G31_n224_2 , 0 , buf_G31_n224_1 );
buf_AQFP buf_G32_splitterfromG32_7_( clk_3 , G32 , 0 , buf_G32_splitterfromG32_7 );
buf_AQFP buf_G32_splitterfromG32_6_( clk_5 , buf_G32_splitterfromG32_7 , 0 , buf_G32_splitterfromG32_6 );
buf_AQFP buf_G32_splitterfromG32_5_( clk_7 , buf_G32_splitterfromG32_6 , 0 , buf_G32_splitterfromG32_5 );
buf_AQFP buf_G32_splitterfromG32_4_( clk_1 , buf_G32_splitterfromG32_5 , 0 , buf_G32_splitterfromG32_4 );
buf_AQFP buf_G32_splitterfromG32_3_( clk_3 , buf_G32_splitterfromG32_4 , 0 , buf_G32_splitterfromG32_3 );
buf_AQFP buf_G32_splitterfromG32_2_( clk_5 , buf_G32_splitterfromG32_3 , 0 , buf_G32_splitterfromG32_2 );
buf_AQFP buf_G32_splitterfromG32_1_( clk_7 , buf_G32_splitterfromG32_2 , 0 , buf_G32_splitterfromG32_1 );
buf_AQFP buf_G33_n260_1_( clk_3 , G33 , 0 , buf_G33_n260_1 );
buf_AQFP buf_G34_n252_1_( clk_3 , G34 , 0 , buf_G34_n252_1 );
buf_AQFP buf_G35_n247_2_( clk_3 , G35 , 0 , buf_G35_n247_2 );
buf_AQFP buf_G35_n247_1_( clk_5 , buf_G35_n247_2 , 0 , buf_G35_n247_1 );
buf_AQFP buf_G36_n199_1_( clk_3 , G36 , 0 , buf_G36_n199_1 );
buf_AQFP buf_G37_n208_1_( clk_3 , G37 , 0 , buf_G37_n208_1 );
buf_AQFP buf_G38_n216_1_( clk_3 , G38 , 0 , buf_G38_n216_1 );
buf_AQFP buf_G39_n238_1_( clk_3 , G39 , 0 , buf_G39_n238_1 );
buf_AQFP buf_G40_n268_1_( clk_3 , G40 , 0 , buf_G40_n268_1 );
buf_AQFP buf_G41_n429_2_( clk_3 , G41 , 0 , buf_G41_n429_2 );
buf_AQFP buf_G41_n429_1_( clk_5 , buf_G41_n429_2 , 0 , buf_G41_n429_1 );
buf_AQFP buf_G42_n228_2_( clk_3 , G42 , 0 , buf_G42_n228_2 );
buf_AQFP buf_G42_n228_1_( clk_5 , buf_G42_n228_2 , 0 , buf_G42_n228_1 );
buf_AQFP buf_G43_splitterfromG43_6_( clk_3 , G43 , 0 , buf_G43_splitterfromG43_6 );
buf_AQFP buf_G43_splitterfromG43_5_( clk_5 , buf_G43_splitterfromG43_6 , 0 , buf_G43_splitterfromG43_5 );
buf_AQFP buf_G43_splitterfromG43_4_( clk_7 , buf_G43_splitterfromG43_5 , 0 , buf_G43_splitterfromG43_4 );
buf_AQFP buf_G43_splitterfromG43_3_( clk_1 , buf_G43_splitterfromG43_4 , 0 , buf_G43_splitterfromG43_3 );
buf_AQFP buf_G43_splitterfromG43_2_( clk_3 , buf_G43_splitterfromG43_3 , 0 , buf_G43_splitterfromG43_2 );
buf_AQFP buf_G43_splitterfromG43_1_( clk_5 , buf_G43_splitterfromG43_2 , 0 , buf_G43_splitterfromG43_1 );
buf_AQFP buf_G44_n264_2_( clk_3 , G44 , 0 , buf_G44_n264_2 );
buf_AQFP buf_G44_n264_1_( clk_5 , buf_G44_n264_2 , 0 , buf_G44_n264_1 );
buf_AQFP buf_G45_n256_2_( clk_3 , G45 , 0 , buf_G45_n256_2 );
buf_AQFP buf_G45_n256_1_( clk_5 , buf_G45_n256_2 , 0 , buf_G45_n256_1 );
buf_AQFP buf_G46_n204_1_( clk_3 , G46 , 0 , buf_G46_n204_1 );
buf_AQFP buf_G47_n212_2_( clk_3 , G47 , 0 , buf_G47_n212_2 );
buf_AQFP buf_G47_n212_1_( clk_5 , buf_G47_n212_2 , 0 , buf_G47_n212_1 );
buf_AQFP buf_G48_n220_2_( clk_3 , G48 , 0 , buf_G48_n220_2 );
buf_AQFP buf_G48_n220_1_( clk_5 , buf_G48_n220_2 , 0 , buf_G48_n220_1 );
buf_AQFP buf_G49_n242_2_( clk_3 , G49 , 0 , buf_G49_n242_2 );
buf_AQFP buf_G49_n242_1_( clk_5 , buf_G49_n242_2 , 0 , buf_G49_n242_1 );
buf_AQFP buf_G5_n320_1_( clk_3 , G5 , 0 , buf_G5_n320_1 );
buf_AQFP buf_G50_n272_2_( clk_3 , G50 , 0 , buf_G50_n272_2 );
buf_AQFP buf_G50_n272_1_( clk_5 , buf_G50_n272_2 , 0 , buf_G50_n272_1 );
buf_AQFP buf_G51_n433_2_( clk_3 , G51 , 0 , buf_G51_n433_2 );
buf_AQFP buf_G51_n433_1_( clk_5 , buf_G51_n433_2 , 0 , buf_G51_n433_1 );
buf_AQFP buf_G52_n229_2_( clk_3 , G52 , 0 , buf_G52_n229_2 );
buf_AQFP buf_G52_n229_1_( clk_5 , buf_G52_n229_2 , 0 , buf_G52_n229_1 );
buf_AQFP buf_G53_splitterfromG53_6_( clk_3 , G53 , 0 , buf_G53_splitterfromG53_6 );
buf_AQFP buf_G53_splitterfromG53_5_( clk_5 , buf_G53_splitterfromG53_6 , 0 , buf_G53_splitterfromG53_5 );
buf_AQFP buf_G53_splitterfromG53_4_( clk_7 , buf_G53_splitterfromG53_5 , 0 , buf_G53_splitterfromG53_4 );
buf_AQFP buf_G53_splitterfromG53_3_( clk_1 , buf_G53_splitterfromG53_4 , 0 , buf_G53_splitterfromG53_3 );
buf_AQFP buf_G53_splitterfromG53_2_( clk_3 , buf_G53_splitterfromG53_3 , 0 , buf_G53_splitterfromG53_2 );
buf_AQFP buf_G53_splitterfromG53_1_( clk_5 , buf_G53_splitterfromG53_2 , 0 , buf_G53_splitterfromG53_1 );
buf_AQFP buf_G54_n265_2_( clk_3 , G54 , 0 , buf_G54_n265_2 );
buf_AQFP buf_G54_n265_1_( clk_5 , buf_G54_n265_2 , 0 , buf_G54_n265_1 );
buf_AQFP buf_G55_n257_2_( clk_3 , G55 , 0 , buf_G55_n257_2 );
buf_AQFP buf_G55_n257_1_( clk_5 , buf_G55_n257_2 , 0 , buf_G55_n257_1 );
buf_AQFP buf_G56_n246_2_( clk_3 , G56 , 0 , buf_G56_n246_2 );
buf_AQFP buf_G56_n246_1_( clk_5 , buf_G56_n246_2 , 0 , buf_G56_n246_1 );
buf_AQFP buf_G57_n205_2_( clk_3 , G57 , 0 , buf_G57_n205_2 );
buf_AQFP buf_G57_n205_1_( clk_5 , buf_G57_n205_2 , 0 , buf_G57_n205_1 );
buf_AQFP buf_G58_n213_2_( clk_3 , G58 , 0 , buf_G58_n213_2 );
buf_AQFP buf_G58_n213_1_( clk_5 , buf_G58_n213_2 , 0 , buf_G58_n213_1 );
buf_AQFP buf_G59_n221_2_( clk_3 , G59 , 0 , buf_G59_n221_2 );
buf_AQFP buf_G59_n221_1_( clk_5 , buf_G59_n221_2 , 0 , buf_G59_n221_1 );
buf_AQFP buf_G6_n404_3_( clk_3 , G6 , 0 , buf_G6_n404_3 );
buf_AQFP buf_G6_n404_2_( clk_5 , buf_G6_n404_3 , 0 , buf_G6_n404_2 );
buf_AQFP buf_G6_n404_1_( clk_7 , buf_G6_n404_2 , 0 , buf_G6_n404_1 );
buf_AQFP buf_G60_n243_2_( clk_3 , G60 , 0 , buf_G60_n243_2 );
buf_AQFP buf_G60_n243_1_( clk_5 , buf_G60_n243_2 , 0 , buf_G60_n243_1 );
buf_AQFP buf_G61_n273_2_( clk_3 , G61 , 0 , buf_G61_n273_2 );
buf_AQFP buf_G61_n273_1_( clk_5 , buf_G61_n273_2 , 0 , buf_G61_n273_1 );
buf_AQFP buf_G62_n434_2_( clk_3 , G62 , 0 , buf_G62_n434_2 );
buf_AQFP buf_G62_n434_1_( clk_5 , buf_G62_n434_2 , 0 , buf_G62_n434_1 );
buf_AQFP buf_G63_n225_1_( clk_3 , G63 , 0 , buf_G63_n225_1 );
buf_AQFP buf_G64_splitterfromG64_6_( clk_3 , G64 , 0 , buf_G64_splitterfromG64_6 );
buf_AQFP buf_G64_splitterfromG64_5_( clk_5 , buf_G64_splitterfromG64_6 , 0 , buf_G64_splitterfromG64_5 );
buf_AQFP buf_G64_splitterfromG64_4_( clk_7 , buf_G64_splitterfromG64_5 , 0 , buf_G64_splitterfromG64_4 );
buf_AQFP buf_G64_splitterfromG64_3_( clk_1 , buf_G64_splitterfromG64_4 , 0 , buf_G64_splitterfromG64_3 );
buf_AQFP buf_G64_splitterfromG64_2_( clk_3 , buf_G64_splitterfromG64_3 , 0 , buf_G64_splitterfromG64_2 );
buf_AQFP buf_G64_splitterfromG64_1_( clk_5 , buf_G64_splitterfromG64_2 , 0 , buf_G64_splitterfromG64_1 );
buf_AQFP buf_G66_n253_1_( clk_3 , G66 , 0 , buf_G66_n253_1 );
buf_AQFP buf_G67_n248_1_( clk_3 , G67 , 0 , buf_G67_n248_1 );
buf_AQFP buf_G68_n200_1_( clk_3 , G68 , 0 , buf_G68_n200_1 );
buf_AQFP buf_G69_n209_1_( clk_3 , G69 , 0 , buf_G69_n209_1 );
buf_AQFP buf_G70_n217_1_( clk_3 , G70 , 0 , buf_G70_n217_1 );
buf_AQFP buf_G71_n239_1_( clk_3 , G71 , 0 , buf_G71_n239_1 );
buf_AQFP buf_G72_n269_1_( clk_3 , G72 , 0 , buf_G72_n269_1 );
buf_AQFP buf_G73_n430_1_( clk_3 , G73 , 0 , buf_G73_n430_1 );
buf_AQFP buf_G74_n163_1_( clk_3 , G74 , 0 , buf_G74_n163_1 );
buf_AQFP buf_G75_n300_2_( clk_3 , G75 , 0 , buf_G75_n300_2 );
buf_AQFP buf_G75_n300_1_( clk_5 , buf_G75_n300_2 , 0 , buf_G75_n300_1 );
buf_AQFP buf_G76_splitterfromG76_6_( clk_3 , G76 , 0 , buf_G76_splitterfromG76_6 );
buf_AQFP buf_G76_splitterfromG76_5_( clk_5 , buf_G76_splitterfromG76_6 , 0 , buf_G76_splitterfromG76_5 );
buf_AQFP buf_G76_splitterfromG76_4_( clk_7 , buf_G76_splitterfromG76_5 , 0 , buf_G76_splitterfromG76_4 );
buf_AQFP buf_G76_splitterfromG76_3_( clk_1 , buf_G76_splitterfromG76_4 , 0 , buf_G76_splitterfromG76_3 );
buf_AQFP buf_G76_splitterfromG76_2_( clk_3 , buf_G76_splitterfromG76_3 , 0 , buf_G76_splitterfromG76_2 );
buf_AQFP buf_G76_splitterfromG76_1_( clk_5 , buf_G76_splitterfromG76_2 , 0 , buf_G76_splitterfromG76_1 );
buf_AQFP buf_G77_n288_2_( clk_3 , G77 , 0 , buf_G77_n288_2 );
buf_AQFP buf_G77_n288_1_( clk_5 , buf_G77_n288_2 , 0 , buf_G77_n288_1 );
buf_AQFP buf_G78_n189_2_( clk_3 , G78 , 0 , buf_G78_n189_2 );
buf_AQFP buf_G78_n189_1_( clk_5 , buf_G78_n189_2 , 0 , buf_G78_n189_1 );
buf_AQFP buf_G79_n179_1_( clk_3 , G79 , 0 , buf_G79_n179_1 );
buf_AQFP buf_G8_splitterG8ton451n486_5_( clk_3 , G8 , 0 , buf_G8_splitterG8ton451n486_5 );
buf_AQFP buf_G8_splitterG8ton451n486_4_( clk_5 , buf_G8_splitterG8ton451n486_5 , 0 , buf_G8_splitterG8ton451n486_4 );
buf_AQFP buf_G8_splitterG8ton451n486_3_( clk_7 , buf_G8_splitterG8ton451n486_4 , 0 , buf_G8_splitterG8ton451n486_3 );
buf_AQFP buf_G8_splitterG8ton451n486_2_( clk_1 , buf_G8_splitterG8ton451n486_3 , 0 , buf_G8_splitterG8ton451n486_2 );
buf_AQFP buf_G8_splitterG8ton451n486_1_( clk_3 , buf_G8_splitterG8ton451n486_2 , 0 , buf_G8_splitterG8ton451n486_1 );
buf_AQFP buf_G80_n192_1_( clk_3 , G80 , 0 , buf_G80_n192_1 );
buf_AQFP buf_G81_n387_2_( clk_3 , G81 , 0 , buf_G81_n387_2 );
buf_AQFP buf_G81_n387_1_( clk_5 , buf_G81_n387_2 , 0 , buf_G81_n387_1 );
buf_AQFP buf_G82_n372_2_( clk_3 , G82 , 0 , buf_G82_n372_2 );
buf_AQFP buf_G82_n372_1_( clk_5 , buf_G82_n372_2 , 0 , buf_G82_n372_1 );
buf_AQFP buf_G83_n357_2_( clk_3 , G83 , 0 , buf_G83_n357_2 );
buf_AQFP buf_G83_n357_1_( clk_5 , buf_G83_n357_2 , 0 , buf_G83_n357_1 );
buf_AQFP buf_G85_n301_2_( clk_3 , G85 , 0 , buf_G85_n301_2 );
buf_AQFP buf_G85_n301_1_( clk_5 , buf_G85_n301_2 , 0 , buf_G85_n301_1 );
buf_AQFP buf_G86_splitterfromG86_7_( clk_3 , G86 , 0 , buf_G86_splitterfromG86_7 );
buf_AQFP buf_G86_splitterfromG86_6_( clk_5 , buf_G86_splitterfromG86_7 , 0 , buf_G86_splitterfromG86_6 );
buf_AQFP buf_G86_splitterfromG86_5_( clk_7 , buf_G86_splitterfromG86_6 , 0 , buf_G86_splitterfromG86_5 );
buf_AQFP buf_G86_splitterfromG86_4_( clk_1 , buf_G86_splitterfromG86_5 , 0 , buf_G86_splitterfromG86_4 );
buf_AQFP buf_G86_splitterfromG86_3_( clk_3 , buf_G86_splitterfromG86_4 , 0 , buf_G86_splitterfromG86_3 );
buf_AQFP buf_G86_splitterfromG86_2_( clk_5 , buf_G86_splitterfromG86_3 , 0 , buf_G86_splitterfromG86_2 );
buf_AQFP buf_G86_splitterfromG86_1_( clk_7 , buf_G86_splitterfromG86_2 , 0 , buf_G86_splitterfromG86_1 );
buf_AQFP buf_G87_n292_2_( clk_3 , G87 , 0 , buf_G87_n292_2 );
buf_AQFP buf_G87_n292_1_( clk_5 , buf_G87_n292_2 , 0 , buf_G87_n292_1 );
buf_AQFP buf_G88_n188_2_( clk_3 , G88 , 0 , buf_G88_n188_2 );
buf_AQFP buf_G88_n188_1_( clk_5 , buf_G88_n188_2 , 0 , buf_G88_n188_1 );
buf_AQFP buf_G89_n181_1_( clk_3 , G89 , 0 , buf_G89_n181_1 );
buf_AQFP buf_G9_n410_1_( clk_3 , G9 , 0 , buf_G9_n410_1 );
buf_AQFP buf_G90_n193_1_( clk_3 , G90 , 0 , buf_G90_n193_1 );
buf_AQFP buf_G91_n391_2_( clk_3 , G91 , 0 , buf_G91_n391_2 );
buf_AQFP buf_G91_n391_1_( clk_5 , buf_G91_n391_2 , 0 , buf_G91_n391_1 );
buf_AQFP buf_G92_n376_2_( clk_3 , G92 , 0 , buf_G92_n376_2 );
buf_AQFP buf_G92_n376_1_( clk_5 , buf_G92_n376_2 , 0 , buf_G92_n376_1 );
buf_AQFP buf_G93_n353_2_( clk_3 , G93 , 0 , buf_G93_n353_2 );
buf_AQFP buf_G93_n353_1_( clk_5 , buf_G93_n353_2 , 0 , buf_G93_n353_1 );
buf_AQFP buf_G95_n303_2_( clk_3 , G95 , 0 , buf_G95_n303_2 );
buf_AQFP buf_G95_n303_1_( clk_5 , buf_G95_n303_2 , 0 , buf_G95_n303_1 );
buf_AQFP buf_G96_splitterfromG96_7_( clk_3 , G96 , 0 , buf_G96_splitterfromG96_7 );
buf_AQFP buf_G96_splitterfromG96_6_( clk_5 , buf_G96_splitterfromG96_7 , 0 , buf_G96_splitterfromG96_6 );
buf_AQFP buf_G96_splitterfromG96_5_( clk_7 , buf_G96_splitterfromG96_6 , 0 , buf_G96_splitterfromG96_5 );
buf_AQFP buf_G96_splitterfromG96_4_( clk_1 , buf_G96_splitterfromG96_5 , 0 , buf_G96_splitterfromG96_4 );
buf_AQFP buf_G96_splitterfromG96_3_( clk_3 , buf_G96_splitterfromG96_4 , 0 , buf_G96_splitterfromG96_3 );
buf_AQFP buf_G96_splitterfromG96_2_( clk_5 , buf_G96_splitterfromG96_3 , 0 , buf_G96_splitterfromG96_2 );
buf_AQFP buf_G96_splitterfromG96_1_( clk_7 , buf_G96_splitterfromG96_2 , 0 , buf_G96_splitterfromG96_1 );
buf_AQFP buf_G97_n289_2_( clk_3 , G97 , 0 , buf_G97_n289_2 );
buf_AQFP buf_G97_n289_1_( clk_5 , buf_G97_n289_2 , 0 , buf_G97_n289_1 );
buf_AQFP buf_G98_n186_2_( clk_3 , G98 , 0 , buf_G98_n186_2 );
buf_AQFP buf_G98_n186_1_( clk_5 , buf_G98_n186_2 , 0 , buf_G98_n186_1 );
buf_AQFP buf_G99_n182_1_( clk_3 , G99 , 0 , buf_G99_n182_1 );
buf_AQFP buf_n160_G2547_8_( clk_7 , n160 , 0 , buf_n160_G2547_8 );
buf_AQFP buf_n160_G2547_7_( clk_1 , buf_n160_G2547_8 , 0 , buf_n160_G2547_7 );
buf_AQFP buf_n160_G2547_6_( clk_3 , buf_n160_G2547_7 , 0 , buf_n160_G2547_6 );
buf_AQFP buf_n160_G2547_5_( clk_5 , buf_n160_G2547_6 , 0 , buf_n160_G2547_5 );
buf_AQFP buf_n160_G2547_4_( clk_7 , buf_n160_G2547_5 , 0 , buf_n160_G2547_4 );
buf_AQFP buf_n160_G2547_3_( clk_1 , buf_n160_G2547_4 , 0 , buf_n160_G2547_3 );
buf_AQFP buf_n160_G2547_2_( clk_3 , buf_n160_G2547_3 , 0 , buf_n160_G2547_2 );
buf_AQFP buf_n160_G2547_1_( clk_5 , buf_n160_G2547_2 , 0 , buf_n160_G2547_1 );
buf_AQFP buf_n162_G2548_12_( clk_6 , n162 , 0 , buf_n162_G2548_12 );
buf_AQFP buf_n162_G2548_11_( clk_8 , buf_n162_G2548_12 , 0 , buf_n162_G2548_11 );
buf_AQFP buf_n162_G2548_10_( clk_2 , buf_n162_G2548_11 , 0 , buf_n162_G2548_10 );
buf_AQFP buf_n162_G2548_9_( clk_4 , buf_n162_G2548_10 , 0 , buf_n162_G2548_9 );
buf_AQFP buf_n162_G2548_8_( clk_6 , buf_n162_G2548_9 , 0 , buf_n162_G2548_8 );
buf_AQFP buf_n162_G2548_7_( clk_8 , buf_n162_G2548_8 , 0 , buf_n162_G2548_7 );
buf_AQFP buf_n162_G2548_6_( clk_2 , buf_n162_G2548_7 , 0 , buf_n162_G2548_6 );
buf_AQFP buf_n162_G2548_5_( clk_4 , buf_n162_G2548_6 , 0 , buf_n162_G2548_5 );
buf_AQFP buf_n162_G2548_4_( clk_6 , buf_n162_G2548_5 , 0 , buf_n162_G2548_4 );
buf_AQFP buf_n162_G2548_3_( clk_8 , buf_n162_G2548_4 , 0 , buf_n162_G2548_3 );
buf_AQFP buf_n162_G2548_2_( clk_2 , buf_n162_G2548_3 , 0 , buf_n162_G2548_2 );
buf_AQFP buf_n162_G2548_1_( clk_4 , buf_n162_G2548_2 , 0 , buf_n162_G2548_1 );
buf_AQFP buf_n163_G2550_12_( clk_6 , n163 , 0 , buf_n163_G2550_12 );
buf_AQFP buf_n163_G2550_11_( clk_8 , buf_n163_G2550_12 , 0 , buf_n163_G2550_11 );
buf_AQFP buf_n163_G2550_10_( clk_2 , buf_n163_G2550_11 , 0 , buf_n163_G2550_10 );
buf_AQFP buf_n163_G2550_9_( clk_4 , buf_n163_G2550_10 , 0 , buf_n163_G2550_9 );
buf_AQFP buf_n163_G2550_8_( clk_6 , buf_n163_G2550_9 , 0 , buf_n163_G2550_8 );
buf_AQFP buf_n163_G2550_7_( clk_8 , buf_n163_G2550_8 , 0 , buf_n163_G2550_7 );
buf_AQFP buf_n163_G2550_6_( clk_2 , buf_n163_G2550_7 , 0 , buf_n163_G2550_6 );
buf_AQFP buf_n163_G2550_5_( clk_4 , buf_n163_G2550_6 , 0 , buf_n163_G2550_5 );
buf_AQFP buf_n163_G2550_4_( clk_6 , buf_n163_G2550_5 , 0 , buf_n163_G2550_4 );
buf_AQFP buf_n163_G2550_3_( clk_8 , buf_n163_G2550_4 , 0 , buf_n163_G2550_3 );
buf_AQFP buf_n163_G2550_2_( clk_2 , buf_n163_G2550_3 , 0 , buf_n163_G2550_2 );
buf_AQFP buf_n163_G2550_1_( clk_4 , buf_n163_G2550_2 , 0 , buf_n163_G2550_1 );
buf_AQFP buf_n164_splittern164ton165G2551_8_( clk_5 , n164 , 0 , buf_n164_splittern164ton165G2551_8 );
buf_AQFP buf_n164_splittern164ton165G2551_7_( clk_7 , buf_n164_splittern164ton165G2551_8 , 0 , buf_n164_splittern164ton165G2551_7 );
buf_AQFP buf_n164_splittern164ton165G2551_6_( clk_1 , buf_n164_splittern164ton165G2551_7 , 0 , buf_n164_splittern164ton165G2551_6 );
buf_AQFP buf_n164_splittern164ton165G2551_5_( clk_3 , buf_n164_splittern164ton165G2551_6 , 0 , buf_n164_splittern164ton165G2551_5 );
buf_AQFP buf_n164_splittern164ton165G2551_4_( clk_5 , buf_n164_splittern164ton165G2551_5 , 0 , buf_n164_splittern164ton165G2551_4 );
buf_AQFP buf_n164_splittern164ton165G2551_3_( clk_7 , buf_n164_splittern164ton165G2551_4 , 0 , buf_n164_splittern164ton165G2551_3 );
buf_AQFP buf_n164_splittern164ton165G2551_2_( clk_1 , buf_n164_splittern164ton165G2551_3 , 0 , buf_n164_splittern164ton165G2551_2 );
buf_AQFP buf_n164_splittern164ton165G2551_1_( clk_3 , buf_n164_splittern164ton165G2551_2 , 0 , buf_n164_splittern164ton165G2551_1 );
buf_AQFP buf_n165_G2552_3_( clk_8 , n165 , 0 , buf_n165_G2552_3 );
buf_AQFP buf_n165_G2552_2_( clk_2 , buf_n165_G2552_3 , 0 , buf_n165_G2552_2 );
buf_AQFP buf_n165_G2552_1_( clk_4 , buf_n165_G2552_2 , 0 , buf_n165_G2552_1 );
buf_AQFP buf_n166_G2553_3_( clk_8 , n166 , 0 , buf_n166_G2553_3 );
buf_AQFP buf_n166_G2553_2_( clk_2 , buf_n166_G2553_3 , 0 , buf_n166_G2553_2 );
buf_AQFP buf_n166_G2553_1_( clk_4 , buf_n166_G2553_2 , 0 , buf_n166_G2553_1 );
buf_AQFP buf_n173_splitterfromn173_2_( clk_1 , n173 , 0 , buf_n173_splitterfromn173_2 );
buf_AQFP buf_n173_splitterfromn173_1_( clk_3 , buf_n173_splitterfromn173_2 , 0 , buf_n173_splitterfromn173_1 );
buf_AQFP buf_n208_n211_1_( clk_6 , n208 , 0 , buf_n208_n211_1 );
buf_AQFP buf_n232_G2563_5_( clk_4 , n232 , 0 , buf_n232_G2563_5 );
buf_AQFP buf_n232_G2563_4_( clk_6 , buf_n232_G2563_5 , 0 , buf_n232_G2563_4 );
buf_AQFP buf_n232_G2563_3_( clk_8 , buf_n232_G2563_4 , 0 , buf_n232_G2563_3 );
buf_AQFP buf_n232_G2563_2_( clk_2 , buf_n232_G2563_3 , 0 , buf_n232_G2563_2 );
buf_AQFP buf_n232_G2563_1_( clk_4 , buf_n232_G2563_2 , 0 , buf_n232_G2563_1 );
buf_AQFP buf_n233_n234_10_( clk_6 , n233 , 0 , buf_n233_n234_10 );
buf_AQFP buf_n233_n234_9_( clk_8 , buf_n233_n234_10 , 0 , buf_n233_n234_9 );
buf_AQFP buf_n233_n234_8_( clk_2 , buf_n233_n234_9 , 0 , buf_n233_n234_8 );
buf_AQFP buf_n233_n234_7_( clk_4 , buf_n233_n234_8 , 0 , buf_n233_n234_7 );
buf_AQFP buf_n233_n234_6_( clk_6 , buf_n233_n234_7 , 0 , buf_n233_n234_6 );
buf_AQFP buf_n233_n234_5_( clk_8 , buf_n233_n234_6 , 0 , buf_n233_n234_5 );
buf_AQFP buf_n233_n234_4_( clk_2 , buf_n233_n234_5 , 0 , buf_n233_n234_4 );
buf_AQFP buf_n233_n234_3_( clk_4 , buf_n233_n234_4 , 0 , buf_n233_n234_3 );
buf_AQFP buf_n233_n234_2_( clk_6 , buf_n233_n234_3 , 0 , buf_n233_n234_2 );
buf_AQFP buf_n233_n234_1_( clk_8 , buf_n233_n234_2 , 0 , buf_n233_n234_1 );
buf_AQFP buf_n236_n237_11_( clk_5 , n236 , 0 , buf_n236_n237_11 );
buf_AQFP buf_n236_n237_10_( clk_7 , buf_n236_n237_11 , 0 , buf_n236_n237_10 );
buf_AQFP buf_n236_n237_9_( clk_1 , buf_n236_n237_10 , 0 , buf_n236_n237_9 );
buf_AQFP buf_n236_n237_8_( clk_3 , buf_n236_n237_9 , 0 , buf_n236_n237_8 );
buf_AQFP buf_n236_n237_7_( clk_5 , buf_n236_n237_8 , 0 , buf_n236_n237_7 );
buf_AQFP buf_n236_n237_6_( clk_7 , buf_n236_n237_7 , 0 , buf_n236_n237_6 );
buf_AQFP buf_n236_n237_5_( clk_1 , buf_n236_n237_6 , 0 , buf_n236_n237_5 );
buf_AQFP buf_n236_n237_4_( clk_3 , buf_n236_n237_5 , 0 , buf_n236_n237_4 );
buf_AQFP buf_n236_n237_3_( clk_5 , buf_n236_n237_4 , 0 , buf_n236_n237_3 );
buf_AQFP buf_n236_n237_2_( clk_7 , buf_n236_n237_3 , 0 , buf_n236_n237_2 );
buf_AQFP buf_n236_n237_1_( clk_1 , buf_n236_n237_2 , 0 , buf_n236_n237_1 );
buf_AQFP buf_n237_G2565_1_( clk_5 , n237 , 0 , buf_n237_G2565_1 );
buf_AQFP buf_n278_splitterfromn278_2_( clk_8 , n278 , 0 , buf_n278_splitterfromn278_2 );
buf_AQFP buf_n278_splitterfromn278_1_( clk_2 , buf_n278_splitterfromn278_2 , 0 , buf_n278_splitterfromn278_1 );
buf_AQFP buf_n281_splitterfromn281_1_( clk_2 , n281 , 0 , buf_n281_splitterfromn281_1 );
buf_AQFP buf_n282_n283_1_( clk_3 , n282 , 0 , buf_n282_n283_1 );
buf_AQFP buf_n283_G2577_4_( clk_6 , n283 , 0 , buf_n283_G2577_4 );
buf_AQFP buf_n283_G2577_3_( clk_8 , buf_n283_G2577_4 , 0 , buf_n283_G2577_3 );
buf_AQFP buf_n283_G2577_2_( clk_2 , buf_n283_G2577_3 , 0 , buf_n283_G2577_2 );
buf_AQFP buf_n283_G2577_1_( clk_4 , buf_n283_G2577_2 , 0 , buf_n283_G2577_1 );
buf_AQFP buf_n287_splitterfromn287_4_( clk_4 , n287 , 0 , buf_n287_splitterfromn287_4 );
buf_AQFP buf_n287_splitterfromn287_3_( clk_6 , buf_n287_splitterfromn287_4 , 0 , buf_n287_splitterfromn287_3 );
buf_AQFP buf_n287_splitterfromn287_2_( clk_8 , buf_n287_splitterfromn287_3 , 0 , buf_n287_splitterfromn287_2 );
buf_AQFP buf_n287_splitterfromn287_1_( clk_2 , buf_n287_splitterfromn287_2 , 0 , buf_n287_splitterfromn287_1 );
buf_AQFP buf_n298_G2580_8_( clk_7 , n298 , 0 , buf_n298_G2580_8 );
buf_AQFP buf_n298_G2580_7_( clk_1 , buf_n298_G2580_8 , 0 , buf_n298_G2580_7 );
buf_AQFP buf_n298_G2580_6_( clk_3 , buf_n298_G2580_7 , 0 , buf_n298_G2580_6 );
buf_AQFP buf_n298_G2580_5_( clk_5 , buf_n298_G2580_6 , 0 , buf_n298_G2580_5 );
buf_AQFP buf_n298_G2580_4_( clk_7 , buf_n298_G2580_5 , 0 , buf_n298_G2580_4 );
buf_AQFP buf_n298_G2580_3_( clk_1 , buf_n298_G2580_4 , 0 , buf_n298_G2580_3 );
buf_AQFP buf_n298_G2580_2_( clk_3 , buf_n298_G2580_3 , 0 , buf_n298_G2580_2 );
buf_AQFP buf_n298_G2580_1_( clk_5 , buf_n298_G2580_2 , 0 , buf_n298_G2580_1 );
buf_AQFP buf_n299_n308_2_( clk_1 , n299 , 0 , buf_n299_n308_2 );
buf_AQFP buf_n299_n308_1_( clk_3 , buf_n299_n308_2 , 0 , buf_n299_n308_1 );
buf_AQFP buf_n310_n312_3_( clk_5 , n310 , 0 , buf_n310_n312_3 );
buf_AQFP buf_n310_n312_2_( clk_7 , buf_n310_n312_3 , 0 , buf_n310_n312_2 );
buf_AQFP buf_n310_n312_1_( clk_1 , buf_n310_n312_2 , 0 , buf_n310_n312_1 );
buf_AQFP buf_n314_n316_2_( clk_7 , n314 , 0 , buf_n314_n316_2 );
buf_AQFP buf_n314_n316_1_( clk_1 , buf_n314_n316_2 , 0 , buf_n314_n316_1 );
buf_AQFP buf_n320_n322_2_( clk_7 , n320 , 0 , buf_n320_n322_2 );
buf_AQFP buf_n320_n322_1_( clk_1 , buf_n320_n322_2 , 0 , buf_n320_n322_1 );
buf_AQFP buf_n324_n326_1_( clk_8 , n324 , 0 , buf_n324_n326_1 );
buf_AQFP buf_n329_n331_2_( clk_8 , n329 , 0 , buf_n329_n331_2 );
buf_AQFP buf_n329_n331_1_( clk_2 , buf_n329_n331_2 , 0 , buf_n329_n331_1 );
buf_AQFP buf_n335_n337_2_( clk_1 , n335 , 0 , buf_n335_n337_2 );
buf_AQFP buf_n335_n337_1_( clk_3 , buf_n335_n337_2 , 0 , buf_n335_n337_1 );
buf_AQFP buf_n339_n341_4_( clk_5 , n339 , 0 , buf_n339_n341_4 );
buf_AQFP buf_n339_n341_3_( clk_7 , buf_n339_n341_4 , 0 , buf_n339_n341_3 );
buf_AQFP buf_n339_n341_2_( clk_1 , buf_n339_n341_3 , 0 , buf_n339_n341_2 );
buf_AQFP buf_n339_n341_1_( clk_3 , buf_n339_n341_2 , 0 , buf_n339_n341_1 );
buf_AQFP buf_n352_n361_3_( clk_6 , n352 , 0 , buf_n352_n361_3 );
buf_AQFP buf_n352_n361_2_( clk_8 , buf_n352_n361_3 , 0 , buf_n352_n361_2 );
buf_AQFP buf_n352_n361_1_( clk_2 , buf_n352_n361_2 , 0 , buf_n352_n361_1 );
buf_AQFP buf_n386_n395_3_( clk_6 , n386 , 0 , buf_n386_n395_3 );
buf_AQFP buf_n386_n395_2_( clk_8 , buf_n386_n395_3 , 0 , buf_n386_n395_2 );
buf_AQFP buf_n386_n395_1_( clk_2 , buf_n386_n395_2 , 0 , buf_n386_n395_1 );
buf_AQFP buf_n398_n400_2_( clk_8 , n398 , 0 , buf_n398_n400_2 );
buf_AQFP buf_n398_n400_1_( clk_2 , buf_n398_n400_2 , 0 , buf_n398_n400_1 );
buf_AQFP buf_n404_n406_1_( clk_2 , n404 , 0 , buf_n404_n406_1 );
buf_AQFP buf_n410_n411_4_( clk_6 , n410 , 0 , buf_n410_n411_4 );
buf_AQFP buf_n410_n411_3_( clk_8 , buf_n410_n411_4 , 0 , buf_n410_n411_3 );
buf_AQFP buf_n410_n411_2_( clk_2 , buf_n410_n411_3 , 0 , buf_n410_n411_2 );
buf_AQFP buf_n410_n411_1_( clk_4 , buf_n410_n411_2 , 0 , buf_n410_n411_1 );
buf_AQFP buf_n420_n422_2_( clk_1 , n420 , 0 , buf_n420_n422_2 );
buf_AQFP buf_n420_n422_1_( clk_3 , buf_n420_n422_2 , 0 , buf_n420_n422_1 );
buf_AQFP buf_n428_splitterfromn428_3_( clk_7 , n428 , 0 , buf_n428_splitterfromn428_3 );
buf_AQFP buf_n428_splitterfromn428_2_( clk_1 , buf_n428_splitterfromn428_3 , 0 , buf_n428_splitterfromn428_2 );
buf_AQFP buf_n428_splitterfromn428_1_( clk_3 , buf_n428_splitterfromn428_2 , 0 , buf_n428_splitterfromn428_1 );
buf_AQFP buf_n436_splitterfromn436_2_( clk_4 , n436 , 0 , buf_n436_splitterfromn436_2 );
buf_AQFP buf_n436_splitterfromn436_1_( clk_6 , buf_n436_splitterfromn436_2 , 0 , buf_n436_splitterfromn436_1 );
buf_AQFP buf_n438_G2586_5_( clk_4 , n438 , 0 , buf_n438_G2586_5 );
buf_AQFP buf_n438_G2586_4_( clk_6 , buf_n438_G2586_5 , 0 , buf_n438_G2586_4 );
buf_AQFP buf_n438_G2586_3_( clk_8 , buf_n438_G2586_4 , 0 , buf_n438_G2586_3 );
buf_AQFP buf_n438_G2586_2_( clk_2 , buf_n438_G2586_3 , 0 , buf_n438_G2586_2 );
buf_AQFP buf_n438_G2586_1_( clk_4 , buf_n438_G2586_2 , 0 , buf_n438_G2586_1 );
buf_AQFP buf_n445_splitterfromn445_4_( clk_3 , n445 , 0 , buf_n445_splitterfromn445_4 );
buf_AQFP buf_n445_splitterfromn445_3_( clk_5 , buf_n445_splitterfromn445_4 , 0 , buf_n445_splitterfromn445_3 );
buf_AQFP buf_n445_splitterfromn445_2_( clk_7 , buf_n445_splitterfromn445_3 , 0 , buf_n445_splitterfromn445_2 );
buf_AQFP buf_n445_splitterfromn445_1_( clk_1 , buf_n445_splitterfromn445_2 , 0 , buf_n445_splitterfromn445_1 );
buf_AQFP buf_n447_splitterfromn447_2_( clk_8 , n447 , 0 , buf_n447_splitterfromn447_2 );
buf_AQFP buf_n447_splitterfromn447_1_( clk_2 , buf_n447_splitterfromn447_2 , 0 , buf_n447_splitterfromn447_1 );
buf_AQFP buf_n452_n498_5_( clk_2 , n452 , 0 , buf_n452_n498_5 );
buf_AQFP buf_n452_n498_4_( clk_4 , buf_n452_n498_5 , 0 , buf_n452_n498_4 );
buf_AQFP buf_n452_n498_3_( clk_6 , buf_n452_n498_4 , 0 , buf_n452_n498_3 );
buf_AQFP buf_n452_n498_2_( clk_8 , buf_n452_n498_3 , 0 , buf_n452_n498_2 );
buf_AQFP buf_n452_n498_1_( clk_2 , buf_n452_n498_2 , 0 , buf_n452_n498_1 );
buf_AQFP buf_n454_n497_2_( clk_6 , n454 , 0 , buf_n454_n497_2 );
buf_AQFP buf_n454_n497_1_( clk_8 , buf_n454_n497_2 , 0 , buf_n454_n497_1 );
buf_AQFP buf_n455_n496_4_( clk_2 , n455 , 0 , buf_n455_n496_4 );
buf_AQFP buf_n455_n496_3_( clk_4 , buf_n455_n496_4 , 0 , buf_n455_n496_3 );
buf_AQFP buf_n455_n496_2_( clk_6 , buf_n455_n496_3 , 0 , buf_n455_n496_2 );
buf_AQFP buf_n455_n496_1_( clk_8 , buf_n455_n496_2 , 0 , buf_n455_n496_1 );
buf_AQFP buf_n517_n518_3_( clk_7 , n517 , 0 , buf_n517_n518_3 );
buf_AQFP buf_n517_n518_2_( clk_1 , buf_n517_n518_3 , 0 , buf_n517_n518_2 );
buf_AQFP buf_n517_n518_1_( clk_3 , buf_n517_n518_2 , 0 , buf_n517_n518_1 );
buf_AQFP buf_n522_n523_3_( clk_7 , n522 , 0 , buf_n522_n523_3 );
buf_AQFP buf_n522_n523_2_( clk_1 , buf_n522_n523_3 , 0 , buf_n522_n523_2 );
buf_AQFP buf_n522_n523_1_( clk_3 , buf_n522_n523_2 , 0 , buf_n522_n523_1 );
buf_AQFP buf_splitterfromG10_G2581_2_( clk_3 , splitterfromG10 , 0 , buf_splitterfromG10_G2581_2 );
buf_AQFP buf_splitterfromG10_G2581_1_( clk_5 , buf_splitterfromG10_G2581_2 , 0 , buf_splitterfromG10_G2581_1 );
buf_AQFP buf_splitterfromG106_G2540_6_( clk_2 , splitterfromG106 , 0 , buf_splitterfromG106_G2540_6 );
buf_AQFP buf_splitterfromG106_G2540_5_( clk_4 , buf_splitterfromG106_G2540_6 , 0 , buf_splitterfromG106_G2540_5 );
buf_AQFP buf_splitterfromG106_G2540_4_( clk_6 , buf_splitterfromG106_G2540_5 , 0 , buf_splitterfromG106_G2540_4 );
buf_AQFP buf_splitterfromG106_G2540_3_( clk_8 , buf_splitterfromG106_G2540_4 , 0 , buf_splitterfromG106_G2540_3 );
buf_AQFP buf_splitterfromG106_G2540_2_( clk_2 , buf_splitterfromG106_G2540_3 , 0 , buf_splitterfromG106_G2540_2 );
buf_AQFP buf_splitterfromG106_G2540_1_( clk_4 , buf_splitterfromG106_G2540_2 , 0 , buf_splitterfromG106_G2540_1 );
buf_AQFP buf_splitterG115ton163G2549_splitterG115toG2531G2549_12_( clk_5 , splitterG115ton163G2549 , 0 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_12 );
buf_AQFP buf_splitterG115ton163G2549_splitterG115toG2531G2549_11_( clk_7 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_12 , 0 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_11 );
buf_AQFP buf_splitterG115ton163G2549_splitterG115toG2531G2549_10_( clk_1 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_11 , 0 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_10 );
buf_AQFP buf_splitterG115ton163G2549_splitterG115toG2531G2549_9_( clk_3 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_10 , 0 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_9 );
buf_AQFP buf_splitterG115ton163G2549_splitterG115toG2531G2549_8_( clk_5 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_9 , 0 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_8 );
buf_AQFP buf_splitterG115ton163G2549_splitterG115toG2531G2549_7_( clk_7 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_8 , 0 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_7 );
buf_AQFP buf_splitterG115ton163G2549_splitterG115toG2531G2549_6_( clk_1 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_7 , 0 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_6 );
buf_AQFP buf_splitterG115ton163G2549_splitterG115toG2531G2549_5_( clk_3 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_6 , 0 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_5 );
buf_AQFP buf_splitterG115ton163G2549_splitterG115toG2531G2549_4_( clk_5 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_5 , 0 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_4 );
buf_AQFP buf_splitterG115ton163G2549_splitterG115toG2531G2549_3_( clk_7 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_4 , 0 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_3 );
buf_AQFP buf_splitterG115ton163G2549_splitterG115toG2531G2549_2_( clk_1 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_3 , 0 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_2 );
buf_AQFP buf_splitterG115ton163G2549_splitterG115toG2531G2549_1_( clk_3 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_2 , 0 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_1 );
buf_AQFP buf_splitterfromG118_n282_1_( clk_7 , splitterfromG118 , 0 , buf_splitterfromG118_n282_1 );
buf_AQFP buf_splitterG123ton284n447_splitterG123ton276n447_1_( clk_8 , splitterG123ton284n447 , 0 , buf_splitterG123ton284n447_splitterG123ton276n447_1 );
buf_AQFP buf_splitterfromG125_n468_1_( clk_6 , splitterfromG125 , 0 , buf_splitterfromG125_n468_1 );
buf_AQFP buf_splitterfromG129_n456_2_( clk_4 , splitterfromG129 , 0 , buf_splitterfromG129_n456_2 );
buf_AQFP buf_splitterfromG129_n456_1_( clk_6 , buf_splitterfromG129_n456_2 , 0 , buf_splitterfromG129_n456_1 );
buf_AQFP buf_splitterfromG130_n480_2_( clk_5 , splitterfromG130 , 0 , buf_splitterfromG130_n480_2 );
buf_AQFP buf_splitterfromG130_n480_1_( clk_7 , buf_splitterfromG130_n480_2 , 0 , buf_splitterfromG130_n480_1 );
buf_AQFP buf_splitterG131ton368n487_n487_1_( clk_6 , splitterG131ton368n487 , 0 , buf_splitterG131ton368n487_n487_1 );
buf_AQFP buf_splitterfromG132_n455_1_( clk_7 , splitterfromG132 , 0 , buf_splitterfromG132_n455_1 );
buf_AQFP buf_splitterfromG133_n452_1_( clk_6 , splitterfromG133 , 0 , buf_splitterfromG133_n452_1 );
buf_AQFP buf_splitterG136ton500n469_splitterG136ton362n469_1_( clk_3 , splitterG136ton500n469 , 0 , buf_splitterG136ton500n469_splitterG136ton362n469_1 );
buf_AQFP buf_splitterG136ton362n469_n469_1_( clk_6 , splitterG136ton362n469 , 0 , buf_splitterG136ton362n469_n469_1 );
buf_AQFP buf_splitterG140ton327n457_n457_1_( clk_5 , splitterG140ton327n457 , 0 , buf_splitterG140ton327n457_n457_1 );
buf_AQFP buf_splitterG141ton158n481_n481_2_( clk_4 , splitterG141ton158n481 , 0 , buf_splitterG141ton158n481_n481_2 );
buf_AQFP buf_splitterG141ton158n481_n481_1_( clk_6 , buf_splitterG141ton158n481_n481_2 , 0 , buf_splitterG141ton158n481_n481_1 );
buf_AQFP buf_splitterG142ton332n488_n488_2_( clk_5 , splitterG142ton332n488 , 0 , buf_splitterG142ton332n488_n488_2 );
buf_AQFP buf_splitterG142ton332n488_n488_1_( clk_7 , buf_splitterG142ton332n488_n488_2 , 0 , buf_splitterG142ton332n488_n488_1 );
buf_AQFP buf_splitterfromG32_G2539_6_( clk_3 , splitterfromG32 , 0 , buf_splitterfromG32_G2539_6 );
buf_AQFP buf_splitterfromG32_G2539_5_( clk_5 , buf_splitterfromG32_G2539_6 , 0 , buf_splitterfromG32_G2539_5 );
buf_AQFP buf_splitterfromG32_G2539_4_( clk_7 , buf_splitterfromG32_G2539_5 , 0 , buf_splitterfromG32_G2539_4 );
buf_AQFP buf_splitterfromG32_G2539_3_( clk_1 , buf_splitterfromG32_G2539_4 , 0 , buf_splitterfromG32_G2539_3 );
buf_AQFP buf_splitterfromG32_G2539_2_( clk_3 , buf_splitterfromG32_G2539_3 , 0 , buf_splitterfromG32_G2539_2 );
buf_AQFP buf_splitterfromG32_G2539_1_( clk_5 , buf_splitterfromG32_G2539_2 , 0 , buf_splitterfromG32_G2539_1 );
buf_AQFP buf_splitterfromG43_G2545_7_( clk_1 , splitterfromG43 , 0 , buf_splitterfromG43_G2545_7 );
buf_AQFP buf_splitterfromG43_G2545_6_( clk_3 , buf_splitterfromG43_G2545_7 , 0 , buf_splitterfromG43_G2545_6 );
buf_AQFP buf_splitterfromG43_G2545_5_( clk_5 , buf_splitterfromG43_G2545_6 , 0 , buf_splitterfromG43_G2545_5 );
buf_AQFP buf_splitterfromG43_G2545_4_( clk_7 , buf_splitterfromG43_G2545_5 , 0 , buf_splitterfromG43_G2545_4 );
buf_AQFP buf_splitterfromG43_G2545_3_( clk_1 , buf_splitterfromG43_G2545_4 , 0 , buf_splitterfromG43_G2545_3 );
buf_AQFP buf_splitterfromG43_G2545_2_( clk_3 , buf_splitterfromG43_G2545_3 , 0 , buf_splitterfromG43_G2545_2 );
buf_AQFP buf_splitterfromG43_G2545_1_( clk_5 , buf_splitterfromG43_G2545_2 , 0 , buf_splitterfromG43_G2545_1 );
buf_AQFP buf_splitterfromG53_G2543_7_( clk_1 , splitterfromG53 , 0 , buf_splitterfromG53_G2543_7 );
buf_AQFP buf_splitterfromG53_G2543_6_( clk_3 , buf_splitterfromG53_G2543_7 , 0 , buf_splitterfromG53_G2543_6 );
buf_AQFP buf_splitterfromG53_G2543_5_( clk_5 , buf_splitterfromG53_G2543_6 , 0 , buf_splitterfromG53_G2543_5 );
buf_AQFP buf_splitterfromG53_G2543_4_( clk_7 , buf_splitterfromG53_G2543_5 , 0 , buf_splitterfromG53_G2543_4 );
buf_AQFP buf_splitterfromG53_G2543_3_( clk_1 , buf_splitterfromG53_G2543_4 , 0 , buf_splitterfromG53_G2543_3 );
buf_AQFP buf_splitterfromG53_G2543_2_( clk_3 , buf_splitterfromG53_G2543_3 , 0 , buf_splitterfromG53_G2543_2 );
buf_AQFP buf_splitterfromG53_G2543_1_( clk_5 , buf_splitterfromG53_G2543_2 , 0 , buf_splitterfromG53_G2543_1 );
buf_AQFP buf_splitterfromG64_G2541_7_( clk_1 , splitterfromG64 , 0 , buf_splitterfromG64_G2541_7 );
buf_AQFP buf_splitterfromG64_G2541_6_( clk_3 , buf_splitterfromG64_G2541_7 , 0 , buf_splitterfromG64_G2541_6 );
buf_AQFP buf_splitterfromG64_G2541_5_( clk_5 , buf_splitterfromG64_G2541_6 , 0 , buf_splitterfromG64_G2541_5 );
buf_AQFP buf_splitterfromG64_G2541_4_( clk_7 , buf_splitterfromG64_G2541_5 , 0 , buf_splitterfromG64_G2541_4 );
buf_AQFP buf_splitterfromG64_G2541_3_( clk_1 , buf_splitterfromG64_G2541_4 , 0 , buf_splitterfromG64_G2541_3 );
buf_AQFP buf_splitterfromG64_G2541_2_( clk_3 , buf_splitterfromG64_G2541_3 , 0 , buf_splitterfromG64_G2541_2 );
buf_AQFP buf_splitterfromG64_G2541_1_( clk_5 , buf_splitterfromG64_G2541_2 , 0 , buf_splitterfromG64_G2541_1 );
buf_AQFP buf_splitterfromG76_G2542_7_( clk_1 , splitterfromG76 , 0 , buf_splitterfromG76_G2542_7 );
buf_AQFP buf_splitterfromG76_G2542_6_( clk_3 , buf_splitterfromG76_G2542_7 , 0 , buf_splitterfromG76_G2542_6 );
buf_AQFP buf_splitterfromG76_G2542_5_( clk_5 , buf_splitterfromG76_G2542_6 , 0 , buf_splitterfromG76_G2542_5 );
buf_AQFP buf_splitterfromG76_G2542_4_( clk_7 , buf_splitterfromG76_G2542_5 , 0 , buf_splitterfromG76_G2542_4 );
buf_AQFP buf_splitterfromG76_G2542_3_( clk_1 , buf_splitterfromG76_G2542_4 , 0 , buf_splitterfromG76_G2542_3 );
buf_AQFP buf_splitterfromG76_G2542_2_( clk_3 , buf_splitterfromG76_G2542_3 , 0 , buf_splitterfromG76_G2542_2 );
buf_AQFP buf_splitterfromG76_G2542_1_( clk_5 , buf_splitterfromG76_G2542_2 , 0 , buf_splitterfromG76_G2542_1 );
buf_AQFP buf_splitterfromG86_G2546_6_( clk_2 , splitterfromG86 , 0 , buf_splitterfromG86_G2546_6 );
buf_AQFP buf_splitterfromG86_G2546_5_( clk_4 , buf_splitterfromG86_G2546_6 , 0 , buf_splitterfromG86_G2546_5 );
buf_AQFP buf_splitterfromG86_G2546_4_( clk_6 , buf_splitterfromG86_G2546_5 , 0 , buf_splitterfromG86_G2546_4 );
buf_AQFP buf_splitterfromG86_G2546_3_( clk_8 , buf_splitterfromG86_G2546_4 , 0 , buf_splitterfromG86_G2546_3 );
buf_AQFP buf_splitterfromG86_G2546_2_( clk_2 , buf_splitterfromG86_G2546_3 , 0 , buf_splitterfromG86_G2546_2 );
buf_AQFP buf_splitterfromG86_G2546_1_( clk_4 , buf_splitterfromG86_G2546_2 , 0 , buf_splitterfromG86_G2546_1 );
buf_AQFP buf_splitterfromG96_G2544_6_( clk_2 , splitterfromG96 , 0 , buf_splitterfromG96_G2544_6 );
buf_AQFP buf_splitterfromG96_G2544_5_( clk_4 , buf_splitterfromG96_G2544_6 , 0 , buf_splitterfromG96_G2544_5 );
buf_AQFP buf_splitterfromG96_G2544_4_( clk_6 , buf_splitterfromG96_G2544_5 , 0 , buf_splitterfromG96_G2544_4 );
buf_AQFP buf_splitterfromG96_G2544_3_( clk_8 , buf_splitterfromG96_G2544_4 , 0 , buf_splitterfromG96_G2544_3 );
buf_AQFP buf_splitterfromG96_G2544_2_( clk_2 , buf_splitterfromG96_G2544_3 , 0 , buf_splitterfromG96_G2544_2 );
buf_AQFP buf_splitterfromG96_G2544_1_( clk_4 , buf_splitterfromG96_G2544_2 , 0 , buf_splitterfromG96_G2544_1 );
buf_AQFP buf_splittern164ton165G2551_G2551_4_( clk_6 , splittern164ton165G2551 , 0 , buf_splittern164ton165G2551_G2551_4 );
buf_AQFP buf_splittern164ton165G2551_G2551_3_( clk_8 , buf_splittern164ton165G2551_G2551_4 , 0 , buf_splittern164ton165G2551_G2551_3 );
buf_AQFP buf_splittern164ton165G2551_G2551_2_( clk_2 , buf_splittern164ton165G2551_G2551_3 , 0 , buf_splittern164ton165G2551_G2551_2 );
buf_AQFP buf_splittern164ton165G2551_G2551_1_( clk_4 , buf_splittern164ton165G2551_G2551_2 , 0 , buf_splittern164ton165G2551_G2551_1 );
buf_AQFP buf_splittern176ton524G2556_G2556_1_( clk_4 , splittern176ton524G2556 , 0 , buf_splittern176ton524G2556_G2556_1 );
buf_AQFP buf_splittern184ton345G2557_splittern184ton442G2557_2_( clk_2 , splittern184ton345G2557 , 0 , buf_splittern184ton345G2557_splittern184ton442G2557_2 );
buf_AQFP buf_splittern184ton345G2557_splittern184ton442G2557_1_( clk_4 , buf_splittern184ton345G2557_splittern184ton442G2557_2 , 0 , buf_splittern184ton345G2557_splittern184ton442G2557_1 );
buf_AQFP buf_splittern184ton442G2557_G2557_8_( clk_7 , splittern184ton442G2557 , 0 , buf_splittern184ton442G2557_G2557_8 );
buf_AQFP buf_splittern184ton442G2557_G2557_7_( clk_1 , buf_splittern184ton442G2557_G2557_8 , 0 , buf_splittern184ton442G2557_G2557_7 );
buf_AQFP buf_splittern184ton442G2557_G2557_6_( clk_3 , buf_splittern184ton442G2557_G2557_7 , 0 , buf_splittern184ton442G2557_G2557_6 );
buf_AQFP buf_splittern184ton442G2557_G2557_5_( clk_5 , buf_splittern184ton442G2557_G2557_6 , 0 , buf_splittern184ton442G2557_G2557_5 );
buf_AQFP buf_splittern184ton442G2557_G2557_4_( clk_7 , buf_splittern184ton442G2557_G2557_5 , 0 , buf_splittern184ton442G2557_G2557_4 );
buf_AQFP buf_splittern184ton442G2557_G2557_3_( clk_1 , buf_splittern184ton442G2557_G2557_4 , 0 , buf_splittern184ton442G2557_G2557_3 );
buf_AQFP buf_splittern184ton442G2557_G2557_2_( clk_3 , buf_splittern184ton442G2557_G2557_3 , 0 , buf_splittern184ton442G2557_G2557_2 );
buf_AQFP buf_splittern184ton442G2557_G2557_1_( clk_5 , buf_splittern184ton442G2557_G2557_2 , 0 , buf_splittern184ton442G2557_G2557_1 );
buf_AQFP buf_splittern191ton330G2558_G2558_9_( clk_4 , splittern191ton330G2558 , 0 , buf_splittern191ton330G2558_G2558_9 );
buf_AQFP buf_splittern191ton330G2558_G2558_8_( clk_6 , buf_splittern191ton330G2558_G2558_9 , 0 , buf_splittern191ton330G2558_G2558_8 );
buf_AQFP buf_splittern191ton330G2558_G2558_7_( clk_8 , buf_splittern191ton330G2558_G2558_8 , 0 , buf_splittern191ton330G2558_G2558_7 );
buf_AQFP buf_splittern191ton330G2558_G2558_6_( clk_2 , buf_splittern191ton330G2558_G2558_7 , 0 , buf_splittern191ton330G2558_G2558_6 );
buf_AQFP buf_splittern191ton330G2558_G2558_5_( clk_4 , buf_splittern191ton330G2558_G2558_6 , 0 , buf_splittern191ton330G2558_G2558_5 );
buf_AQFP buf_splittern191ton330G2558_G2558_4_( clk_6 , buf_splittern191ton330G2558_G2558_5 , 0 , buf_splittern191ton330G2558_G2558_4 );
buf_AQFP buf_splittern191ton330G2558_G2558_3_( clk_8 , buf_splittern191ton330G2558_G2558_4 , 0 , buf_splittern191ton330G2558_G2558_3 );
buf_AQFP buf_splittern191ton330G2558_G2558_2_( clk_2 , buf_splittern191ton330G2558_G2558_3 , 0 , buf_splittern191ton330G2558_G2558_2 );
buf_AQFP buf_splittern191ton330G2558_G2558_1_( clk_4 , buf_splittern191ton330G2558_G2558_2 , 0 , buf_splittern191ton330G2558_G2558_1 );
buf_AQFP buf_splittern198ton325G2559_G2559_10_( clk_2 , splittern198ton325G2559 , 0 , buf_splittern198ton325G2559_G2559_10 );
buf_AQFP buf_splittern198ton325G2559_G2559_9_( clk_4 , buf_splittern198ton325G2559_G2559_10 , 0 , buf_splittern198ton325G2559_G2559_9 );
buf_AQFP buf_splittern198ton325G2559_G2559_8_( clk_6 , buf_splittern198ton325G2559_G2559_9 , 0 , buf_splittern198ton325G2559_G2559_8 );
buf_AQFP buf_splittern198ton325G2559_G2559_7_( clk_8 , buf_splittern198ton325G2559_G2559_8 , 0 , buf_splittern198ton325G2559_G2559_7 );
buf_AQFP buf_splittern198ton325G2559_G2559_6_( clk_2 , buf_splittern198ton325G2559_G2559_7 , 0 , buf_splittern198ton325G2559_G2559_6 );
buf_AQFP buf_splittern198ton325G2559_G2559_5_( clk_4 , buf_splittern198ton325G2559_G2559_6 , 0 , buf_splittern198ton325G2559_G2559_5 );
buf_AQFP buf_splittern198ton325G2559_G2559_4_( clk_6 , buf_splittern198ton325G2559_G2559_5 , 0 , buf_splittern198ton325G2559_G2559_4 );
buf_AQFP buf_splittern198ton325G2559_G2559_3_( clk_8 , buf_splittern198ton325G2559_G2559_4 , 0 , buf_splittern198ton325G2559_G2559_3 );
buf_AQFP buf_splittern198ton325G2559_G2559_2_( clk_2 , buf_splittern198ton325G2559_G2559_3 , 0 , buf_splittern198ton325G2559_G2559_2 );
buf_AQFP buf_splittern198ton325G2559_G2559_1_( clk_4 , buf_splittern198ton325G2559_G2559_2 , 0 , buf_splittern198ton325G2559_G2559_1 );
buf_AQFP buf_splittern207ton366G2569_splittern207ton486G2569_2_( clk_3 , splittern207ton366G2569 , 0 , buf_splittern207ton366G2569_splittern207ton486G2569_2 );
buf_AQFP buf_splittern207ton366G2569_splittern207ton486G2569_1_( clk_5 , buf_splittern207ton366G2569_splittern207ton486G2569_2 , 0 , buf_splittern207ton366G2569_splittern207ton486G2569_1 );
buf_AQFP buf_splittern207ton486G2569_splittern207toG2560G2569_6_( clk_8 , splittern207ton486G2569 , 0 , buf_splittern207ton486G2569_splittern207toG2560G2569_6 );
buf_AQFP buf_splittern207ton486G2569_splittern207toG2560G2569_5_( clk_2 , buf_splittern207ton486G2569_splittern207toG2560G2569_6 , 0 , buf_splittern207ton486G2569_splittern207toG2560G2569_5 );
buf_AQFP buf_splittern207ton486G2569_splittern207toG2560G2569_4_( clk_4 , buf_splittern207ton486G2569_splittern207toG2560G2569_5 , 0 , buf_splittern207ton486G2569_splittern207toG2560G2569_4 );
buf_AQFP buf_splittern207ton486G2569_splittern207toG2560G2569_3_( clk_6 , buf_splittern207ton486G2569_splittern207toG2560G2569_4 , 0 , buf_splittern207ton486G2569_splittern207toG2560G2569_3 );
buf_AQFP buf_splittern207ton486G2569_splittern207toG2560G2569_2_( clk_8 , buf_splittern207ton486G2569_splittern207toG2560G2569_3 , 0 , buf_splittern207ton486G2569_splittern207toG2560G2569_2 );
buf_AQFP buf_splittern207ton486G2569_splittern207toG2560G2569_1_( clk_2 , buf_splittern207ton486G2569_splittern207toG2560G2569_2 , 0 , buf_splittern207ton486G2569_splittern207toG2560G2569_1 );
buf_AQFP buf_splittern215ton315G2568_splittern215ton479G2568_2_( clk_3 , splittern215ton315G2568 , 0 , buf_splittern215ton315G2568_splittern215ton479G2568_2 );
buf_AQFP buf_splittern215ton315G2568_splittern215ton479G2568_1_( clk_5 , buf_splittern215ton315G2568_splittern215ton479G2568_2 , 0 , buf_splittern215ton315G2568_splittern215ton479G2568_1 );
buf_AQFP buf_splittern215ton479G2568_splittern215ton280G2568_2_( clk_8 , splittern215ton479G2568 , 0 , buf_splittern215ton479G2568_splittern215ton280G2568_2 );
buf_AQFP buf_splittern215ton479G2568_splittern215ton280G2568_1_( clk_2 , buf_splittern215ton479G2568_splittern215ton280G2568_2 , 0 , buf_splittern215ton479G2568_splittern215ton280G2568_1 );
buf_AQFP buf_splittern215ton280G2568_splittern215toG2561G2568_3_( clk_6 , splittern215ton280G2568 , 0 , buf_splittern215ton280G2568_splittern215toG2561G2568_3 );
buf_AQFP buf_splittern215ton280G2568_splittern215toG2561G2568_2_( clk_8 , buf_splittern215ton280G2568_splittern215toG2561G2568_3 , 0 , buf_splittern215ton280G2568_splittern215toG2561G2568_2 );
buf_AQFP buf_splittern215ton280G2568_splittern215toG2561G2568_1_( clk_2 , buf_splittern215ton280G2568_splittern215toG2561G2568_2 , 0 , buf_splittern215ton280G2568_splittern215toG2561G2568_1 );
buf_AQFP buf_splittern223ton321G2567_splittern223ton459G2567_3_( clk_3 , splittern223ton321G2567 , 0 , buf_splittern223ton321G2567_splittern223ton459G2567_3 );
buf_AQFP buf_splittern223ton321G2567_splittern223ton459G2567_2_( clk_5 , buf_splittern223ton321G2567_splittern223ton459G2567_3 , 0 , buf_splittern223ton321G2567_splittern223ton459G2567_2 );
buf_AQFP buf_splittern223ton321G2567_splittern223ton459G2567_1_( clk_7 , buf_splittern223ton321G2567_splittern223ton459G2567_2 , 0 , buf_splittern223ton321G2567_splittern223ton459G2567_1 );
buf_AQFP buf_splittern223ton277G2567_splittern223toG2562G2567_4_( clk_4 , splittern223ton277G2567 , 0 , buf_splittern223ton277G2567_splittern223toG2562G2567_4 );
buf_AQFP buf_splittern223ton277G2567_splittern223toG2562G2567_3_( clk_6 , buf_splittern223ton277G2567_splittern223toG2562G2567_4 , 0 , buf_splittern223ton277G2567_splittern223toG2562G2567_3 );
buf_AQFP buf_splittern223ton277G2567_splittern223toG2562G2567_2_( clk_8 , buf_splittern223ton277G2567_splittern223toG2562G2567_3 , 0 , buf_splittern223ton277G2567_splittern223toG2562G2567_2 );
buf_AQFP buf_splittern223ton277G2567_splittern223toG2562G2567_1_( clk_2 , buf_splittern223ton277G2567_splittern223toG2562G2567_2 , 0 , buf_splittern223ton277G2567_splittern223toG2562G2567_1 );
buf_AQFP buf_splittern231ton311n232_splittern231ton284n232_2_( clk_3 , splittern231ton311n232 , 0 , buf_splittern231ton311n232_splittern231ton284n232_2 );
buf_AQFP buf_splittern231ton311n232_splittern231ton284n232_1_( clk_5 , buf_splittern231ton311n232_splittern231ton284n232_2 , 0 , buf_splittern231ton311n232_splittern231ton284n232_1 );
buf_AQFP buf_splittern245ton336G2566_splittern245ton474G2566_2_( clk_4 , splittern245ton336G2566 , 0 , buf_splittern245ton336G2566_splittern245ton474G2566_2 );
buf_AQFP buf_splittern245ton336G2566_splittern245ton474G2566_1_( clk_6 , buf_splittern245ton336G2566_splittern245ton474G2566_2 , 0 , buf_splittern245ton336G2566_splittern245ton474G2566_1 );
buf_AQFP buf_splittern245ton474G2566_splittern245ton279G2566_1_( clk_2 , splittern245ton474G2566 , 0 , buf_splittern245ton474G2566_splittern245ton279G2566_1 );
buf_AQFP buf_splittern245ton279G2566_G2566_4_( clk_6 , splittern245ton279G2566 , 0 , buf_splittern245ton279G2566_G2566_4 );
buf_AQFP buf_splittern245ton279G2566_G2566_3_( clk_8 , buf_splittern245ton279G2566_G2566_4 , 0 , buf_splittern245ton279G2566_G2566_3 );
buf_AQFP buf_splittern245ton279G2566_G2566_2_( clk_2 , buf_splittern245ton279G2566_G2566_3 , 0 , buf_splittern245ton279G2566_G2566_2 );
buf_AQFP buf_splittern245ton279G2566_G2566_1_( clk_4 , buf_splittern245ton279G2566_G2566_2 , 0 , buf_splittern245ton279G2566_G2566_1 );
buf_AQFP buf_splittern251ton421G2570_splittern251ton493G2570_4_( clk_4 , splittern251ton421G2570 , 0 , buf_splittern251ton421G2570_splittern251ton493G2570_4 );
buf_AQFP buf_splittern251ton421G2570_splittern251ton493G2570_3_( clk_6 , buf_splittern251ton421G2570_splittern251ton493G2570_4 , 0 , buf_splittern251ton421G2570_splittern251ton493G2570_3 );
buf_AQFP buf_splittern251ton421G2570_splittern251ton493G2570_2_( clk_8 , buf_splittern251ton421G2570_splittern251ton493G2570_3 , 0 , buf_splittern251ton421G2570_splittern251ton493G2570_2 );
buf_AQFP buf_splittern251ton421G2570_splittern251ton493G2570_1_( clk_2 , buf_splittern251ton421G2570_splittern251ton493G2570_2 , 0 , buf_splittern251ton421G2570_splittern251ton493G2570_1 );
buf_AQFP buf_splittern251ton493G2570_G2570_5_( clk_5 , splittern251ton493G2570 , 0 , buf_splittern251ton493G2570_G2570_5 );
buf_AQFP buf_splittern251ton493G2570_G2570_4_( clk_7 , buf_splittern251ton493G2570_G2570_5 , 0 , buf_splittern251ton493G2570_G2570_4 );
buf_AQFP buf_splittern251ton493G2570_G2570_3_( clk_1 , buf_splittern251ton493G2570_G2570_4 , 0 , buf_splittern251ton493G2570_G2570_3 );
buf_AQFP buf_splittern251ton493G2570_G2570_2_( clk_3 , buf_splittern251ton493G2570_G2570_3 , 0 , buf_splittern251ton493G2570_G2570_2 );
buf_AQFP buf_splittern251ton493G2570_G2570_1_( clk_5 , buf_splittern251ton493G2570_G2570_2 , 0 , buf_splittern251ton493G2570_G2570_1 );
buf_AQFP buf_splittern259ton405G2571_splittern259ton454G2571_4_( clk_4 , splittern259ton405G2571 , 0 , buf_splittern259ton405G2571_splittern259ton454G2571_4 );
buf_AQFP buf_splittern259ton405G2571_splittern259ton454G2571_3_( clk_6 , buf_splittern259ton405G2571_splittern259ton454G2571_4 , 0 , buf_splittern259ton405G2571_splittern259ton454G2571_3 );
buf_AQFP buf_splittern259ton405G2571_splittern259ton454G2571_2_( clk_8 , buf_splittern259ton405G2571_splittern259ton454G2571_3 , 0 , buf_splittern259ton405G2571_splittern259ton454G2571_2 );
buf_AQFP buf_splittern259ton405G2571_splittern259ton454G2571_1_( clk_2 , buf_splittern259ton405G2571_splittern259ton454G2571_2 , 0 , buf_splittern259ton405G2571_splittern259ton454G2571_1 );
buf_AQFP buf_splittern259ton454G2571_G2571_5_( clk_5 , splittern259ton454G2571 , 0 , buf_splittern259ton454G2571_G2571_5 );
buf_AQFP buf_splittern259ton454G2571_G2571_4_( clk_7 , buf_splittern259ton454G2571_G2571_5 , 0 , buf_splittern259ton454G2571_G2571_4 );
buf_AQFP buf_splittern259ton454G2571_G2571_3_( clk_1 , buf_splittern259ton454G2571_G2571_4 , 0 , buf_splittern259ton454G2571_G2571_3 );
buf_AQFP buf_splittern259ton454G2571_G2571_2_( clk_3 , buf_splittern259ton454G2571_G2571_3 , 0 , buf_splittern259ton454G2571_G2571_2 );
buf_AQFP buf_splittern259ton454G2571_G2571_1_( clk_5 , buf_splittern259ton454G2571_G2571_2 , 0 , buf_splittern259ton454G2571_G2571_1 );
buf_AQFP buf_splittern267ton399G2572_G2572_9_( clk_4 , splittern267ton399G2572 , 0 , buf_splittern267ton399G2572_G2572_9 );
buf_AQFP buf_splittern267ton399G2572_G2572_8_( clk_6 , buf_splittern267ton399G2572_G2572_9 , 0 , buf_splittern267ton399G2572_G2572_8 );
buf_AQFP buf_splittern267ton399G2572_G2572_7_( clk_8 , buf_splittern267ton399G2572_G2572_8 , 0 , buf_splittern267ton399G2572_G2572_7 );
buf_AQFP buf_splittern267ton399G2572_G2572_6_( clk_2 , buf_splittern267ton399G2572_G2572_7 , 0 , buf_splittern267ton399G2572_G2572_6 );
buf_AQFP buf_splittern267ton399G2572_G2572_5_( clk_4 , buf_splittern267ton399G2572_G2572_6 , 0 , buf_splittern267ton399G2572_G2572_5 );
buf_AQFP buf_splittern267ton399G2572_G2572_4_( clk_6 , buf_splittern267ton399G2572_G2572_5 , 0 , buf_splittern267ton399G2572_G2572_4 );
buf_AQFP buf_splittern267ton399G2572_G2572_3_( clk_8 , buf_splittern267ton399G2572_G2572_4 , 0 , buf_splittern267ton399G2572_G2572_3 );
buf_AQFP buf_splittern267ton399G2572_G2572_2_( clk_2 , buf_splittern267ton399G2572_G2572_3 , 0 , buf_splittern267ton399G2572_G2572_2 );
buf_AQFP buf_splittern267ton399G2572_G2572_1_( clk_4 , buf_splittern267ton399G2572_G2572_2 , 0 , buf_splittern267ton399G2572_G2572_1 );
buf_AQFP buf_splittern275ton340n283_splittern275ton286n283_1_( clk_4 , splittern275ton340n283 , 0 , buf_splittern275ton340n283_splittern275ton286n283_1 );
buf_AQFP buf_splitterfromn436_n446_2_( clk_1 , splitterfromn436 , 0 , buf_splitterfromn436_n446_2 );
buf_AQFP buf_splitterfromn436_n446_1_( clk_3 , buf_splitterfromn436_n446_2 , 0 , buf_splitterfromn436_n446_1 );
buf_AQFP buf_splitterfromn445_G2587_1_( clk_5 , splitterfromn445 , 0 , buf_splitterfromn445_G2587_1 );
buf_AQFP buf_splittern453ton481n454_splittern453ton493n454_1_( clk_1 , splittern453ton481n454 , 0 , buf_splittern453ton481n454_splittern453ton493n454_1 );
buf_AQFP buf_splittern503ton504n522_n522_2_( clk_2 , splittern503ton504n522 , 0 , buf_splittern503ton504n522_n522_2 );
buf_AQFP buf_splittern503ton504n522_n522_1_( clk_4 , buf_splittern503ton504n522_n522_2 , 0 , buf_splittern503ton504n522_n522_1 );
buf_AQFP buf_splitterfromn505_n519_1_( clk_7 , splitterfromn505 , 0 , buf_splitterfromn505_n519_1 );
splitter_AQFP splitterfromG10_( clk_1 , buf_G10_splitterfromG10_1 , 0 , splitterfromG10 );
splitter_AQFP splitterfromG106_( clk_8 , buf_G106_splitterfromG106_1 , 0 , splitterfromG106 );
splitter_AQFP splitterG115ton163G2549_( clk_3 , G115 , 0 , splitterG115ton163G2549 );
splitter_AQFP splitterG115toG2531G2549_( clk_4 , buf_splitterG115ton163G2549_splitterG115toG2531G2549_1 , 0 , splitterG115toG2531G2549 );
splitter_AQFP splitterG117ton203n429_( clk_2 , G117 , 0 , splitterG117ton203n429 );
splitter_AQFP splitterG117ton199n217_( clk_3 , splitterG117ton203n429 , 0 , splitterG117ton199n217 );
splitter_AQFP splitterG117ton269n429_( clk_3 , splitterG117ton203n429 , 0 , splitterG117ton269n429 );
splitter_AQFP splitterG117ton209n238_( clk_4 , splitterG117ton269n429 , 0 , splitterG117ton209n238 );
splitter_AQFP splitterG117ton239n253_( clk_4 , splitterG117ton269n429 , 0 , splitterG117ton239n253 );
splitter_AQFP splitterG117ton260n429_( clk_4 , splitterG117ton269n429 , 0 , splitterG117ton260n429 );
splitter_AQFP splitterG117ton224n429_( clk_5 , splitterG117ton260n429 , 0 , splitterG117ton224n429 );
splitter_AQFP splitterfromG118_( clk_5 , buf_G118_splitterfromG118_1 , 0 , splitterfromG118 );
splitter_AQFP splitterfromG119_( clk_4 , buf_G119_splitterfromG119_1 , 0 , splitterfromG119 );
splitter_AQFP splitterG12ton310n421_( clk_2 , G12 , 0 , splitterG12ton310n421 );
splitter_AQFP splitterG12ton314n421_( clk_4 , splitterG12ton310n421 , 0 , splitterG12ton314n421 );
splitter_AQFP splitterG12ton335n421_( clk_6 , splitterG12ton314n421 , 0 , splitterG12ton335n421 );
splitter_AQFP splitterG12ton365n421_( clk_8 , splitterG12ton335n421 , 0 , splitterG12ton365n421 );
splitter_AQFP splitterG12ton321n421_( clk_1 , splitterG12ton365n421 , 0 , splitterG12ton321n421 );
splitter_AQFP splitterG12ton340n421_( clk_2 , splitterG12ton321n421 , 0 , splitterG12ton340n421 );
splitter_AQFP splitterG120ton203n431_( clk_2 , G120 , 0 , splitterG120ton203n431 );
splitter_AQFP splitterG120ton262n431_( clk_3 , splitterG120ton203n431 , 0 , splitterG120ton262n431 );
splitter_AQFP splitterG120ton270n431_( clk_4 , splitterG120ton262n431 , 0 , splitterG120ton270n431 );
splitter_AQFP splitterG120ton240n431_( clk_5 , splitterG120ton270n431 , 0 , splitterG120ton240n431 );
splitter_AQFP splitterG121ton161n233_( clk_2 , G121 , 0 , splitterG121ton161n233 );
splitter_AQFP splitterG122ton437n438_( clk_6 , buf_G122_splitterG122ton437n438_1 , 0 , splitterG122ton437n438 );
splitter_AQFP splitterG122ton282n438_( clk_8 , splitterG122ton437n438 , 0 , splitterG122ton282n438 );
splitter_AQFP splitterG123ton285n447_( clk_4 , buf_G123_splitterG123ton285n447_1 , 0 , splitterG123ton285n447 );
splitter_AQFP splitterG123ton284n447_( clk_6 , splitterG123ton285n447 , 0 , splitterG123ton284n447 );
splitter_AQFP splitterG123ton276n447_( clk_2 , buf_splitterG123ton284n447_splitterG123ton276n447_1 , 0 , splitterG123ton276n447 );
splitter_AQFP splitterG123ton446n447_( clk_4 , splitterG123ton276n447 , 0 , splitterG123ton446n447 );
splitter_AQFP splitterfromG124_( clk_4 , buf_G124_splitterfromG124_1 , 0 , splitterfromG124 );
splitter_AQFP splitterfromG125_( clk_4 , buf_G125_splitterfromG125_1 , 0 , splitterfromG125 );
splitter_AQFP splitterfromG126_( clk_3 , buf_G126_splitterfromG126_1 , 0 , splitterfromG126 );
splitter_AQFP splitterfromG128_( clk_3 , buf_G128_splitterfromG128_1 , 0 , splitterfromG128 );
splitter_AQFP splitterfromG129_( clk_2 , buf_G129_splitterfromG129_1 , 0 , splitterfromG129 );
splitter_AQFP splitterfromG130_( clk_3 , buf_G130_splitterfromG130_1 , 0 , splitterfromG130 );
splitter_AQFP splitterG131ton368n487_( clk_4 , buf_G131_splitterG131ton368n487_1 , 0 , splitterG131ton368n487 );
splitter_AQFP splitterfromG132_( clk_5 , buf_G132_splitterfromG132_1 , 0 , splitterfromG132 );
splitter_AQFP splitterfromG133_( clk_4 , buf_G133_splitterfromG133_1 , 0 , splitterfromG133 );
splitter_AQFP splitterG134ton513n401_( clk_1 , buf_G134_splitterG134ton513n401_1 , 0 , splitterG134ton513n401 );
splitter_AQFP splitterG134ton506n401_( clk_3 , splitterG134ton513n401 , 0 , splitterG134ton506n401 );
splitter_AQFP splitterG135ton505n309_( clk_1 , buf_G135_splitterG135ton505n309_1 , 0 , splitterG135ton505n309 );
splitter_AQFP splitterG135ton510n309_( clk_3 , splitterG135ton505n309 , 0 , splitterG135ton510n309 );
splitter_AQFP splitterG136ton500n469_( clk_1 , buf_G136_splitterG136ton500n469_1 , 0 , splitterG136ton500n469 );
splitter_AQFP splitterG136ton362n469_( clk_4 , buf_splitterG136ton500n469_splitterG136ton362n469_1 , 0 , splitterG136ton362n469 );
splitter_AQFP splitterG137toG2536G2538_( clk_4 , buf_G137_splitterG137toG2536G2538_1 , 0 , splitterG137toG2536G2538 );
splitter_AQFP splitterG138ton502n465_( clk_2 , buf_G138_splitterG138ton502n465_1 , 0 , splitterG138ton502n465 );
splitter_AQFP splitterG138ton381n465_( clk_4 , splitterG138ton502n465 , 0 , splitterG138ton381n465 );
splitter_AQFP splitterG139ton159n461_( clk_1 , buf_G139_splitterG139ton159n461_1 , 0 , splitterG139ton159n461 );
splitter_AQFP splitterG139ton396n461_( clk_3 , splitterG139ton159n461 , 0 , splitterG139ton396n461 );
splitter_AQFP splitterG140ton159n457_( clk_1 , buf_G140_splitterG140ton159n457_1 , 0 , splitterG140ton159n457 );
splitter_AQFP splitterG140ton327n457_( clk_3 , splitterG140ton159n457 , 0 , splitterG140ton327n457 );
splitter_AQFP splitterG141ton158n481_( clk_2 , buf_G141_splitterG141ton158n481_1 , 0 , splitterG141ton158n481 );
splitter_AQFP splitterG142ton158n488_( clk_1 , buf_G142_splitterG142ton158n488_1 , 0 , splitterG142ton158n488 );
splitter_AQFP splitterG142ton332n488_( clk_3 , splitterG142ton158n488 , 0 , splitterG142ton332n488 );
splitter_AQFP splitterfromG143_( clk_1 , buf_G143_splitterfromG143_1 , 0 , splitterfromG143 );
splitter_AQFP splitterfromG147_( clk_4 , buf_G147_splitterfromG147_1 , 0 , splitterfromG147 );
splitter_AQFP splitterG23ton409n408_( clk_2 , G23 , 0 , splitterG23ton409n408 );
splitter_AQFP splitterG23ton352n408_( clk_3 , splitterG23ton409n408 , 0 , splitterG23ton352n408 );
splitter_AQFP splitterG23ton299n408_( clk_5 , splitterG23ton352n408 , 0 , splitterG23ton299n408 );
splitter_AQFP splitterG23ton344n408_( clk_7 , splitterG23ton299n408 , 0 , splitterG23ton344n408 );
splitter_AQFP splitterG23ton371n408_( clk_1 , splitterG23ton344n408 , 0 , splitterG23ton371n408 );
splitter_AQFP splitterG23ton330n408_( clk_2 , splitterG23ton371n408 , 0 , splitterG23ton330n408 );
splitter_AQFP splitterfromG32_( clk_1 , buf_G32_splitterfromG32_1 , 0 , splitterfromG32 );
splitter_AQFP splitterfromG43_( clk_7 , buf_G43_splitterfromG43_1 , 0 , splitterfromG43 );
splitter_AQFP splitterfromG53_( clk_7 , buf_G53_splitterfromG53_1 , 0 , splitterfromG53 );
splitter_AQFP splitterfromG64_( clk_7 , buf_G64_splitterfromG64_1 , 0 , splitterfromG64 );
splitter_AQFP splitterfromG76_( clk_7 , buf_G76_splitterfromG76_1 , 0 , splitterfromG76 );
splitter_AQFP splitterG8ton451n486_( clk_4 , buf_G8_splitterG8ton451n486_1 , 0 , splitterG8ton451n486 );
splitter_AQFP splitterG8ton479n486_( clk_6 , splitterG8ton451n486 , 0 , splitterG8ton479n486 );
splitter_AQFP splitterfromG86_( clk_8 , buf_G86_splitterfromG86_1 , 0 , splitterfromG86 );
splitter_AQFP splitterfromG96_( clk_8 , buf_G96_splitterfromG96_1 , 0 , splitterfromG96 );
splitter_AQFP splittern164ton165G2551_( clk_4 , buf_n164_splittern164ton165G2551_1 , 0 , splittern164ton165G2551 );
splitter_AQFP splitterfromn169_( clk_5 , n169 , 0 , splitterfromn169 );
splitter_AQFP splitterfromn172_( clk_5 , n172 , 0 , splitterfromn172 );
splitter_AQFP splitterfromn173_( clk_4 , buf_n173_splitterfromn173_1 , 0 , splitterfromn173 );
splitter_AQFP splittern176ton234G2556_( clk_8 , n176 , 0 , splittern176ton234G2556 );
splitter_AQFP splittern176ton524G2556_( clk_2 , splittern176ton234G2556 , 0 , splittern176ton524G2556 );
splitter_AQFP splittern177ton178n391_( clk_3 , n177 , 0 , splittern177ton178n391 );
splitter_AQFP splittern177ton181n193_( clk_4 , splittern177ton178n391 , 0 , splittern177ton181n193 );
splitter_AQFP splittern177ton195n391_( clk_4 , splittern177ton178n391 , 0 , splittern177ton195n391 );
splitter_AQFP splittern177ton373n291_( clk_5 , splittern177ton195n391 , 0 , splittern177ton373n291 );
splitter_AQFP splittern177ton185n188_( clk_6 , splittern177ton373n291 , 0 , splittern177ton185n188 );
splitter_AQFP splittern177ton189n291_( clk_6 , splittern177ton373n291 , 0 , splittern177ton189n291 );
splitter_AQFP splittern177ton292n391_( clk_5 , splittern177ton195n391 , 0 , splittern177ton292n391 );
splitter_AQFP splittern177ton292n303_( clk_6 , splittern177ton292n391 , 0 , splittern177ton292n303 );
splitter_AQFP splittern177ton304n356_( clk_6 , splittern177ton292n391 , 0 , splittern177ton304n356 );
splitter_AQFP splittern177ton357n376_( clk_6 , splittern177ton292n391 , 0 , splittern177ton357n376 );
splitter_AQFP splittern177ton387n391_( clk_6 , splittern177ton292n391 , 0 , splittern177ton387n391 );
splitter_AQFP splittern184ton345G2557_( clk_8 , n184 , 0 , splittern184ton345G2557 );
splitter_AQFP splittern184ton442G2557_( clk_5 , buf_splittern184ton345G2557_splittern184ton442G2557_1 , 0 , splittern184ton442G2557 );
splitter_AQFP splittern191ton330G2558_( clk_2 , n191 , 0 , splittern191ton330G2558 );
splitter_AQFP splittern198ton325G2559_( clk_8 , n198 , 0 , splittern198ton325G2559 );
splitter_AQFP splittern203ton204n434_( clk_4 , n203 , 0 , splittern203ton204n434 );
splitter_AQFP splittern203ton205n220_( clk_5 , splittern203ton204n434 , 0 , splittern203ton205n220 );
splitter_AQFP splittern203ton221n246_( clk_5 , splittern203ton204n434 , 0 , splittern203ton221n246 );
splitter_AQFP splittern203ton264n434_( clk_5 , splittern203ton204n434 , 0 , splittern203ton264n434 );
splitter_AQFP splittern203ton242n257_( clk_6 , splittern203ton264n434 , 0 , splittern203ton242n257 );
splitter_AQFP splittern203ton272n434_( clk_6 , splittern203ton264n434 , 0 , splittern203ton272n434 );
splitter_AQFP splittern207ton366G2569_( clk_1 , n207 , 0 , splittern207ton366G2569 );
splitter_AQFP splittern207ton486G2569_( clk_6 , buf_splittern207ton366G2569_splittern207ton486G2569_1 , 0 , splittern207ton486G2569 );
splitter_AQFP splittern207toG2560G2569_( clk_4 , buf_splittern207ton486G2569_splittern207toG2560G2569_1 , 0 , splittern207toG2560G2569 );
splitter_AQFP splittern215ton315G2568_( clk_1 , n215 , 0 , splittern215ton315G2568 );
splitter_AQFP splittern215ton479G2568_( clk_6 , buf_splittern215ton315G2568_splittern215ton479G2568_1 , 0 , splittern215ton479G2568 );
splitter_AQFP splittern215ton280G2568_( clk_4 , buf_splittern215ton479G2568_splittern215ton280G2568_1 , 0 , splittern215ton280G2568 );
splitter_AQFP splittern215toG2561G2568_( clk_4 , buf_splittern215ton280G2568_splittern215toG2561G2568_1 , 0 , splittern215toG2561G2568 );
splitter_AQFP splittern223ton321G2567_( clk_1 , n223 , 0 , splittern223ton321G2567 );
splitter_AQFP splittern223ton459G2567_( clk_8 , buf_splittern223ton321G2567_splittern223ton459G2567_1 , 0 , splittern223ton459G2567 );
splitter_AQFP splittern223ton277G2567_( clk_2 , splittern223ton459G2567 , 0 , splittern223ton277G2567 );
splitter_AQFP splittern223toG2562G2567_( clk_4 , buf_splittern223ton277G2567_splittern223toG2562G2567_1 , 0 , splittern223toG2562G2567 );
splitter_AQFP splittern231ton311n232_( clk_1 , n231 , 0 , splittern231ton311n232 );
splitter_AQFP splittern231ton284n232_( clk_6 , buf_splittern231ton311n232_splittern231ton284n232_1 , 0 , splittern231ton284n232 );
splitter_AQFP splittern231ton471n232_( clk_8 , splittern231ton284n232 , 0 , splittern231ton471n232 );
splitter_AQFP splitterfromn234_( clk_2 , n234 , 0 , splitterfromn234 );
splitter_AQFP splittern245ton336G2566_( clk_2 , n245 , 0 , splittern245ton336G2566 );
splitter_AQFP splittern245ton474G2566_( clk_8 , buf_splittern245ton336G2566_splittern245ton474G2566_1 , 0 , splittern245ton474G2566 );
splitter_AQFP splittern245ton279G2566_( clk_4 , buf_splittern245ton474G2566_splittern245ton279G2566_1 , 0 , splittern245ton279G2566 );
splitter_AQFP splittern251ton421G2570_( clk_2 , n251 , 0 , splittern251ton421G2570 );
splitter_AQFP splittern251ton493G2570_( clk_3 , buf_splittern251ton421G2570_splittern251ton493G2570_1 , 0 , splittern251ton493G2570 );
splitter_AQFP splittern259ton405G2571_( clk_2 , n259 , 0 , splittern259ton405G2571 );
splitter_AQFP splittern259ton454G2571_( clk_3 , buf_splittern259ton405G2571_splittern259ton454G2571_1 , 0 , splittern259ton454G2571 );
splitter_AQFP splittern267ton399G2572_( clk_2 , n267 , 0 , splittern267ton399G2572 );
splitter_AQFP splittern275ton340n283_( clk_2 , n275 , 0 , splittern275ton340n283 );
splitter_AQFP splittern275ton286n283_( clk_6 , buf_splittern275ton340n283_splittern275ton286n283_1 , 0 , splittern275ton286n283 );
splitter_AQFP splittern275ton467n283_( clk_8 , splittern275ton286n283 , 0 , splittern275ton467n283 );
splitter_AQFP splittern275ton276n283_( clk_2 , splittern275ton467n283 , 0 , splittern275ton276n283 );
splitter_AQFP splitterfromn278_( clk_4 , buf_n278_splitterfromn278_1 , 0 , splitterfromn278 );
splitter_AQFP splitterfromn281_( clk_4 , buf_n281_splitterfromn281_1 , 0 , splitterfromn281 );
splitter_AQFP splitterfromn287_( clk_4 , buf_n287_splitterfromn287_1 , 0 , splitterfromn287 );
splitter_AQFP splittern294ton295n440_( clk_2 , n294 , 0 , splittern294ton295n440 );
splitter_AQFP splittern294ton408n440_( clk_3 , splittern294ton295n440 , 0 , splittern294ton408n440 );
splitter_AQFP splittern306ton307n510_( clk_2 , n306 , 0 , splittern306ton307n510 );
splitter_AQFP splitterfromn309_( clk_7 , n309 , 0 , splitterfromn309 );
splitter_AQFP splitterfromn313_( clk_6 , n313 , 0 , splitterfromn313 );
splitter_AQFP splitterfromn317_( clk_5 , n317 , 0 , splitterfromn317 );
splitter_AQFP splitterfromn323_( clk_5 , n323 , 0 , splitterfromn323 );
splitter_AQFP splitterfromn327_( clk_5 , n327 , 0 , splitterfromn327 );
splitter_AQFP splitterfromn332_( clk_6 , n332 , 0 , splitterfromn332 );
splitter_AQFP splitterfromn338_( clk_6 , n338 , 0 , splitterfromn338 );
splitter_AQFP splitterfromn342_( clk_6 , n342 , 0 , splitterfromn342 );
splitter_AQFP splitterfromn347_( clk_4 , n347 , 0 , splitterfromn347 );
splitter_AQFP splitterfromn359_( clk_2 , n359 , 0 , splitterfromn359 );
splitter_AQFP splitterfromn361_( clk_5 , n361 , 0 , splitterfromn361 );
splitter_AQFP splitterfromn367_( clk_4 , n367 , 0 , splitterfromn367 );
splitter_AQFP splitterfromn378_( clk_2 , n378 , 0 , splitterfromn378 );
splitter_AQFP splitterfromn380_( clk_5 , n380 , 0 , splitterfromn380 );
splitter_AQFP splitterfromn396_( clk_5 , n396 , 0 , splitterfromn396 );
splitter_AQFP splitterfromn401_( clk_6 , n401 , 0 , splitterfromn401 );
splitter_AQFP splitterfromn407_( clk_6 , n407 , 0 , splitterfromn407 );
splitter_AQFP splitterfromn428_( clk_4 , buf_n428_splitterfromn428_1 , 0 , splitterfromn428 );
splitter_AQFP splitterfromn436_( clk_7 , buf_n436_splitterfromn436_1 , 0 , splitterfromn436 );
splitter_AQFP splitterfromn441_( clk_6 , n441 , 0 , splitterfromn441 );
splitter_AQFP splitterfromn445_( clk_3 , buf_n445_splitterfromn445_1 , 0 , splitterfromn445 );
splitter_AQFP splitterfromn447_( clk_4 , buf_n447_splitterfromn447_1 , 0 , splitterfromn447 );
splitter_AQFP splitterfromn448_( clk_2 , n448 , 0 , splitterfromn448 );
splitter_AQFP splitterfromn449_( clk_2 , n449 , 0 , splitterfromn449 );
splitter_AQFP splittern450ton460n469_( clk_4 , n450 , 0 , splittern450ton460n469 );
splitter_AQFP splittern450ton451n469_( clk_5 , splittern450ton460n469 , 0 , splittern450ton451n469 );
splitter_AQFP splittern450ton456n469_( clk_6 , splittern450ton451n469 , 0 , splittern450ton456n469 );
splitter_AQFP splittern451ton452n487_( clk_7 , n451 , 0 , splittern451ton452n487 );
splitter_AQFP splittern453ton481n454_( clk_7 , n453 , 0 , splittern453ton481n454 );
splitter_AQFP splittern453ton493n454_( clk_2 , buf_splittern453ton481n454_splittern453ton493n454_1 , 0 , splittern453ton493n454 );
splitter_AQFP splitterfromn459_( clk_3 , n459 , 0 , splitterfromn459 );
splitter_AQFP splitterfromn462_( clk_8 , n462 , 0 , splitterfromn462 );
splitter_AQFP splitterfromn466_( clk_8 , n466 , 0 , splitterfromn466 );
splitter_AQFP splitterfromn483_( clk_3 , n483 , 0 , splitterfromn483 );
splitter_AQFP splitterfromn490_( clk_4 , n490 , 0 , splitterfromn490 );
splitter_AQFP splittern499ton514n512_( clk_4 , n499 , 0 , splittern499ton514n512 );
splitter_AQFP splittern499ton503n512_( clk_5 , splittern499ton514n512 , 0 , splittern499ton503n512 );
splitter_AQFP splitterfromn500_( clk_5 , n500 , 0 , splitterfromn500 );
splitter_AQFP splittern503ton504n522_( clk_8 , n503 , 0 , splittern503ton504n522 );
splitter_AQFP splitterfromn504_( clk_3 , n504 , 0 , splitterfromn504 );
splitter_AQFP splitterfromn505_( clk_5 , n505 , 0 , splitterfromn505 );
splitter_AQFP splitterfromn512_( clk_8 , n512 , 0 , splitterfromn512 );
splitter_AQFP splitterfromn514_( clk_7 , n514 , 0 , splitterfromn514 );
splitter_AQFP splitterfromn525_( clk_5 , n525 , 0 , splitterfromn525 );

endmodule