module top( clk_1 , clk_2 , clk_3 , clk_4 , clk_5 , clk_6 , clk_7 , clk_8 , G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G4 , G5 , G6 , G7 , G8 , G9 , G1884 , G1885 , G1886 , G1887 , G1888 , G1889 , G1890 , G1891 , G1892 , G1893 , G1894 , G1895 , G1896 , G1897 , G1898 , G1899 , G1900 , G1901 , G1902 , G1903 , G1904 , G1905 , G1906 , G1907 , G1908 );

input G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G4 , G5 , G6 , G7 , G8 , G9 ;
output G1884 , G1885 , G1886 , G1887 , G1888 , G1889 , G1890 , G1891 , G1892 , G1893 , G1894 , G1895 , G1896 , G1897 , G1898 , G1899 , G1900 , G1901 , G1902 , G1903 , G1904 , G1905 , G1906 , G1907 , G1908 ;
wire n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , buf_G1_splitterG1ton48n208_1 , buf_G12_splitterG12ton163n259_1 , buf_G16_splitterG16ton64n230_1 , buf_G17_splitterfromG17_1 , buf_G18_splitterfromG18_1 , buf_G19_splitterfromG19_1 , buf_G20_splitterfromG20_1 , buf_G21_splitterfromG21_1 , buf_G22_splitterfromG22_1 , buf_G25_splitterG25ton193n281_8 , buf_G25_splitterG25ton193n281_7 , buf_G25_splitterG25ton193n281_6 , buf_G25_splitterG25ton193n281_5 , buf_G25_splitterG25ton193n281_4 , buf_G25_splitterG25ton193n281_3 , buf_G25_splitterG25ton193n281_2 , buf_G25_splitterG25ton193n281_1 , buf_G26_splitterG26ton100n320_7 , buf_G26_splitterG26ton100n320_6 , buf_G26_splitterG26ton100n320_5 , buf_G26_splitterG26ton100n320_4 , buf_G26_splitterG26ton100n320_3 , buf_G26_splitterG26ton100n320_2 , buf_G26_splitterG26ton100n320_1 , buf_G27_splitterG27ton153n287_7 , buf_G27_splitterG27ton153n287_6 , buf_G27_splitterG27ton153n287_5 , buf_G27_splitterG27ton153n287_4 , buf_G27_splitterG27ton153n287_3 , buf_G27_splitterG27ton153n287_2 , buf_G27_splitterG27ton153n287_1 , buf_G28_splitterG28ton173n291_7 , buf_G28_splitterG28ton173n291_6 , buf_G28_splitterG28ton173n291_5 , buf_G28_splitterG28ton173n291_4 , buf_G28_splitterG28ton173n291_3 , buf_G28_splitterG28ton173n291_2 , buf_G28_splitterG28ton173n291_1 , buf_G29_splitterfromG29_1 , buf_G30_splitterfromG30_1 , buf_G31_splitterG31ton127n282_1 , buf_G32_splitterfromG32_6 , buf_G32_splitterfromG32_5 , buf_G32_splitterfromG32_4 , buf_G32_splitterfromG32_3 , buf_G32_splitterfromG32_2 , buf_G32_splitterfromG32_1 , buf_G5_splitterG5ton143n237_1 , buf_n35_splittern35ton269n252_5 , buf_n35_splittern35ton269n252_4 , buf_n35_splittern35ton269n252_3 , buf_n35_splittern35ton269n252_2 , buf_n35_splittern35ton269n252_1 , buf_n74_splittern74ton75n275_5 , buf_n74_splittern74ton75n275_4 , buf_n74_splittern74ton75n275_3 , buf_n74_splittern74ton75n275_2 , buf_n74_splittern74ton75n275_1 , buf_n128_splittern128ton129n295_4 , buf_n128_splittern128ton129n295_3 , buf_n128_splittern128ton129n295_2 , buf_n128_splittern128ton129n295_1 , buf_n178_splittern178ton269n232_5 , buf_n178_splittern178ton269n232_4 , buf_n178_splittern178ton269n232_3 , buf_n178_splittern178ton269n232_2 , buf_n178_splittern178ton269n232_1 , buf_n199_splitterfromn199_3 , buf_n199_splitterfromn199_2 , buf_n199_splitterfromn199_1 , buf_n200_splitterfromn200_4 , buf_n200_splitterfromn200_3 , buf_n200_splitterfromn200_2 , buf_n200_splitterfromn200_1 , buf_n205_splitterfromn205_1 , buf_n209_G1884_1 , buf_n212_G1885_1 , buf_n215_G1886_1 , buf_n218_G1887_1 , buf_n219_splitterfromn219_2 , buf_n219_splitterfromn219_1 , buf_n221_splittern221ton222n254_1 , buf_n225_G1888_1 , buf_n228_G1889_1 , buf_n231_G1890_1 , buf_n238_G1891_2 , buf_n238_G1891_1 , buf_n241_G1892_1 , buf_n244_G1893_1 , buf_n247_G1894_1 , buf_n251_G1895_2 , buf_n251_G1895_1 , buf_n257_G1896_1 , buf_n260_G1897_1 , buf_n263_G1898_1 , buf_n266_G1899_1 , buf_n272_n273_2 , buf_n272_n273_1 , buf_n274_G1900_1 , buf_n287_n288_5 , buf_n287_n288_4 , buf_n287_n288_3 , buf_n287_n288_2 , buf_n287_n288_1 , buf_n291_n292_4 , buf_n291_n292_3 , buf_n291_n292_2 , buf_n291_n292_1 , buf_n295_n296_4 , buf_n295_n296_3 , buf_n295_n296_2 , buf_n295_n296_1 , buf_n299_splitterfromn299_7 , buf_n299_splitterfromn299_6 , buf_n299_splitterfromn299_5 , buf_n299_splitterfromn299_4 , buf_n299_splitterfromn299_3 , buf_n299_splitterfromn299_2 , buf_n299_splitterfromn299_1 , buf_n300_splitterfromn300_10 , buf_n300_splitterfromn300_9 , buf_n300_splitterfromn300_8 , buf_n300_splitterfromn300_7 , buf_n300_splitterfromn300_6 , buf_n300_splitterfromn300_5 , buf_n300_splitterfromn300_4 , buf_n300_splitterfromn300_3 , buf_n300_splitterfromn300_2 , buf_n300_splitterfromn300_1 , buf_n311_splitterfromn311_7 , buf_n311_splitterfromn311_6 , buf_n311_splitterfromn311_5 , buf_n311_splitterfromn311_4 , buf_n311_splitterfromn311_3 , buf_n311_splitterfromn311_2 , buf_n311_splitterfromn311_1 , buf_n312_splitterfromn312_10 , buf_n312_splitterfromn312_9 , buf_n312_splitterfromn312_8 , buf_n312_splitterfromn312_7 , buf_n312_splitterfromn312_6 , buf_n312_splitterfromn312_5 , buf_n312_splitterfromn312_4 , buf_n312_splitterfromn312_3 , buf_n312_splitterfromn312_2 , buf_n312_splitterfromn312_1 , buf_n321_n322_1 , buf_n322_G1908_1 , buf_splitterG1ton48n208_n48_1 , buf_splitterG1ton49n208_splitterG1ton207n208_11 , buf_splitterG1ton49n208_splitterG1ton207n208_10 , buf_splitterG1ton49n208_splitterG1ton207n208_9 , buf_splitterG1ton49n208_splitterG1ton207n208_8 , buf_splitterG1ton49n208_splitterG1ton207n208_7 , buf_splitterG1ton49n208_splitterG1ton207n208_6 , buf_splitterG1ton49n208_splitterG1ton207n208_5 , buf_splitterG1ton49n208_splitterG1ton207n208_4 , buf_splitterG1ton49n208_splitterG1ton207n208_3 , buf_splitterG1ton49n208_splitterG1ton207n208_2 , buf_splitterG1ton49n208_splitterG1ton207n208_1 , buf_splitterG10ton61n224_splitterG10ton120n224_2 , buf_splitterG10ton61n224_splitterG10ton120n224_1 , buf_splitterG10ton120n224_splitterG10ton223n224_10 , buf_splitterG10ton120n224_splitterG10ton223n224_9 , buf_splitterG10ton120n224_splitterG10ton223n224_8 , buf_splitterG10ton120n224_splitterG10ton223n224_7 , buf_splitterG10ton120n224_splitterG10ton223n224_6 , buf_splitterG10ton120n224_splitterG10ton223n224_5 , buf_splitterG10ton120n224_splitterG10ton223n224_4 , buf_splitterG10ton120n224_splitterG10ton223n224_3 , buf_splitterG10ton120n224_splitterG10ton223n224_2 , buf_splitterG10ton120n224_splitterG10ton223n224_1 , buf_splitterG11ton135n256_splitterG11ton255n256_12 , buf_splitterG11ton135n256_splitterG11ton255n256_11 , buf_splitterG11ton135n256_splitterG11ton255n256_10 , buf_splitterG11ton135n256_splitterG11ton255n256_9 , buf_splitterG11ton135n256_splitterG11ton255n256_8 , buf_splitterG11ton135n256_splitterG11ton255n256_7 , buf_splitterG11ton135n256_splitterG11ton255n256_6 , buf_splitterG11ton135n256_splitterG11ton255n256_5 , buf_splitterG11ton135n256_splitterG11ton255n256_4 , buf_splitterG11ton135n256_splitterG11ton255n256_3 , buf_splitterG11ton135n256_splitterG11ton255n256_2 , buf_splitterG11ton135n256_splitterG11ton255n256_1 , buf_splitterG12ton163n259_n163_1 , buf_splitterG12ton164n259_splitterG12ton258n259_11 , buf_splitterG12ton164n259_splitterG12ton258n259_10 , buf_splitterG12ton164n259_splitterG12ton258n259_9 , buf_splitterG12ton164n259_splitterG12ton258n259_8 , buf_splitterG12ton164n259_splitterG12ton258n259_7 , buf_splitterG12ton164n259_splitterG12ton258n259_6 , buf_splitterG12ton164n259_splitterG12ton258n259_5 , buf_splitterG12ton164n259_splitterG12ton258n259_4 , buf_splitterG12ton164n259_splitterG12ton258n259_3 , buf_splitterG12ton164n259_splitterG12ton258n259_2 , buf_splitterG12ton164n259_splitterG12ton258n259_1 , buf_splitterG13ton79n262_splitterG13ton111n262_1 , buf_splitterG13ton111n262_splitterG13ton261n262_11 , buf_splitterG13ton111n262_splitterG13ton261n262_10 , buf_splitterG13ton111n262_splitterG13ton261n262_9 , buf_splitterG13ton111n262_splitterG13ton261n262_8 , buf_splitterG13ton111n262_splitterG13ton261n262_7 , buf_splitterG13ton111n262_splitterG13ton261n262_6 , buf_splitterG13ton111n262_splitterG13ton261n262_5 , buf_splitterG13ton111n262_splitterG13ton261n262_4 , buf_splitterG13ton111n262_splitterG13ton261n262_3 , buf_splitterG13ton111n262_splitterG13ton261n262_2 , buf_splitterG13ton111n262_splitterG13ton261n262_1 , buf_splitterG14ton103n265_splitterG14ton264n265_12 , buf_splitterG14ton103n265_splitterG14ton264n265_11 , buf_splitterG14ton103n265_splitterG14ton264n265_10 , buf_splitterG14ton103n265_splitterG14ton264n265_9 , buf_splitterG14ton103n265_splitterG14ton264n265_8 , buf_splitterG14ton103n265_splitterG14ton264n265_7 , buf_splitterG14ton103n265_splitterG14ton264n265_6 , buf_splitterG14ton103n265_splitterG14ton264n265_5 , buf_splitterG14ton103n265_splitterG14ton264n265_4 , buf_splitterG14ton103n265_splitterG14ton264n265_3 , buf_splitterG14ton103n265_splitterG14ton264n265_2 , buf_splitterG14ton103n265_splitterG14ton264n265_1 , buf_splitterG15ton135n227_splitterG15ton226n227_13 , buf_splitterG15ton135n227_splitterG15ton226n227_12 , buf_splitterG15ton135n227_splitterG15ton226n227_11 , buf_splitterG15ton135n227_splitterG15ton226n227_10 , buf_splitterG15ton135n227_splitterG15ton226n227_9 , buf_splitterG15ton135n227_splitterG15ton226n227_8 , buf_splitterG15ton135n227_splitterG15ton226n227_7 , buf_splitterG15ton135n227_splitterG15ton226n227_6 , buf_splitterG15ton135n227_splitterG15ton226n227_5 , buf_splitterG15ton135n227_splitterG15ton226n227_4 , buf_splitterG15ton135n227_splitterG15ton226n227_3 , buf_splitterG15ton135n227_splitterG15ton226n227_2 , buf_splitterG15ton135n227_splitterG15ton226n227_1 , buf_splitterG16ton64n230_n64_1 , buf_splitterG16ton65n230_splitterG16ton229n230_11 , buf_splitterG16ton65n230_splitterG16ton229n230_10 , buf_splitterG16ton65n230_splitterG16ton229n230_9 , buf_splitterG16ton65n230_splitterG16ton229n230_8 , buf_splitterG16ton65n230_splitterG16ton229n230_7 , buf_splitterG16ton65n230_splitterG16ton229n230_6 , buf_splitterG16ton65n230_splitterG16ton229n230_5 , buf_splitterG16ton65n230_splitterG16ton229n230_4 , buf_splitterG16ton65n230_splitterG16ton229n230_3 , buf_splitterG16ton65n230_splitterG16ton229n230_2 , buf_splitterG16ton65n230_splitterG16ton229n230_1 , buf_splitterfromG17_n74_1 , buf_splitterfromG18_n35_1 , buf_splitterfromG19_n128_1 , buf_splitterG2ton45n211_splitterG2ton146n211_2 , buf_splitterG2ton45n211_splitterG2ton146n211_1 , buf_splitterG2ton146n211_splitterG2ton210n211_10 , buf_splitterG2ton146n211_splitterG2ton210n211_9 , buf_splitterG2ton146n211_splitterG2ton210n211_8 , buf_splitterG2ton146n211_splitterG2ton210n211_7 , buf_splitterG2ton146n211_splitterG2ton210n211_6 , buf_splitterG2ton146n211_splitterG2ton210n211_5 , buf_splitterG2ton146n211_splitterG2ton210n211_4 , buf_splitterG2ton146n211_splitterG2ton210n211_3 , buf_splitterG2ton146n211_splitterG2ton210n211_2 , buf_splitterG2ton146n211_splitterG2ton210n211_1 , buf_splitterfromG20_n178_1 , buf_splitterG25ton193n281_n281_6 , buf_splitterG25ton193n281_n281_5 , buf_splitterG25ton193n281_n281_4 , buf_splitterG25ton193n281_n281_3 , buf_splitterG25ton193n281_n281_2 , buf_splitterG25ton193n281_n281_1 , buf_splitterG26ton100n320_n320_7 , buf_splitterG26ton100n320_n320_6 , buf_splitterG26ton100n320_n320_5 , buf_splitterG26ton100n320_n320_4 , buf_splitterG26ton100n320_n320_3 , buf_splitterG26ton100n320_n320_2 , buf_splitterG26ton100n320_n320_1 , buf_splitterG27ton153n287_n287_1 , buf_splitterG28ton173n291_n291_2 , buf_splitterG28ton173n291_n291_1 , buf_splitterfromG29_n199_1 , buf_splitterG3ton156n214_splitterG3ton213n214_12 , buf_splitterG3ton156n214_splitterG3ton213n214_11 , buf_splitterG3ton156n214_splitterG3ton213n214_10 , buf_splitterG3ton156n214_splitterG3ton213n214_9 , buf_splitterG3ton156n214_splitterG3ton213n214_8 , buf_splitterG3ton156n214_splitterG3ton213n214_7 , buf_splitterG3ton156n214_splitterG3ton213n214_6 , buf_splitterG3ton156n214_splitterG3ton213n214_5 , buf_splitterG3ton156n214_splitterG3ton213n214_4 , buf_splitterG3ton156n214_splitterG3ton213n214_3 , buf_splitterG3ton156n214_splitterG3ton213n214_2 , buf_splitterG3ton156n214_splitterG3ton213n214_1 , buf_splitterfromG30_n219_1 , buf_splitterG31ton127n282_splitterG31ton126n282_5 , buf_splitterG31ton127n282_splitterG31ton126n282_4 , buf_splitterG31ton127n282_splitterG31ton126n282_3 , buf_splitterG31ton127n282_splitterG31ton126n282_2 , buf_splitterG31ton127n282_splitterG31ton126n282_1 , buf_splitterG31ton291n282_splitterG31ton276n282_4 , buf_splitterG31ton291n282_splitterG31ton276n282_3 , buf_splitterG31ton291n282_splitterG31ton276n282_2 , buf_splitterG31ton291n282_splitterG31ton276n282_1 , buf_splitterfromG32_n268_9 , buf_splitterfromG32_n268_8 , buf_splitterfromG32_n268_7 , buf_splitterfromG32_n268_6 , buf_splitterfromG32_n268_5 , buf_splitterfromG32_n268_4 , buf_splitterfromG32_n268_3 , buf_splitterfromG32_n268_2 , buf_splitterfromG32_n268_1 , buf_splitterG33ton199n316_splitterG33ton203n316_3 , buf_splitterG33ton199n316_splitterG33ton203n316_2 , buf_splitterG33ton199n316_splitterG33ton203n316_1 , buf_splitterG33ton203n316_splitterG33ton273n316_7 , buf_splitterG33ton203n316_splitterG33ton273n316_6 , buf_splitterG33ton203n316_splitterG33ton273n316_5 , buf_splitterG33ton203n316_splitterG33ton273n316_4 , buf_splitterG33ton203n316_splitterG33ton273n316_3 , buf_splitterG33ton203n316_splitterG33ton273n316_2 , buf_splitterG33ton203n316_splitterG33ton273n316_1 , buf_splitterG4ton118n217_splitterG4ton216n217_11 , buf_splitterG4ton118n217_splitterG4ton216n217_10 , buf_splitterG4ton118n217_splitterG4ton216n217_9 , buf_splitterG4ton118n217_splitterG4ton216n217_8 , buf_splitterG4ton118n217_splitterG4ton216n217_7 , buf_splitterG4ton118n217_splitterG4ton216n217_6 , buf_splitterG4ton118n217_splitterG4ton216n217_5 , buf_splitterG4ton118n217_splitterG4ton216n217_4 , buf_splitterG4ton118n217_splitterG4ton216n217_3 , buf_splitterG4ton118n217_splitterG4ton216n217_2 , buf_splitterG4ton118n217_splitterG4ton216n217_1 , buf_splitterG5ton39n237_splitterG5ton236n237_10 , buf_splitterG5ton39n237_splitterG5ton236n237_9 , buf_splitterG5ton39n237_splitterG5ton236n237_8 , buf_splitterG5ton39n237_splitterG5ton236n237_7 , buf_splitterG5ton39n237_splitterG5ton236n237_6 , buf_splitterG5ton39n237_splitterG5ton236n237_5 , buf_splitterG5ton39n237_splitterG5ton236n237_4 , buf_splitterG5ton39n237_splitterG5ton236n237_3 , buf_splitterG5ton39n237_splitterG5ton236n237_2 , buf_splitterG5ton39n237_splitterG5ton236n237_1 , buf_splitterG6ton156n240_splitterG6ton239n240_11 , buf_splitterG6ton156n240_splitterG6ton239n240_10 , buf_splitterG6ton156n240_splitterG6ton239n240_9 , buf_splitterG6ton156n240_splitterG6ton239n240_8 , buf_splitterG6ton156n240_splitterG6ton239n240_7 , buf_splitterG6ton156n240_splitterG6ton239n240_6 , buf_splitterG6ton156n240_splitterG6ton239n240_5 , buf_splitterG6ton156n240_splitterG6ton239n240_4 , buf_splitterG6ton156n240_splitterG6ton239n240_3 , buf_splitterG6ton156n240_splitterG6ton239n240_2 , buf_splitterG6ton156n240_splitterG6ton239n240_1 , buf_splitterG7ton117n243_splitterG7ton242n243_11 , buf_splitterG7ton117n243_splitterG7ton242n243_10 , buf_splitterG7ton117n243_splitterG7ton242n243_9 , buf_splitterG7ton117n243_splitterG7ton242n243_8 , buf_splitterG7ton117n243_splitterG7ton242n243_7 , buf_splitterG7ton117n243_splitterG7ton242n243_6 , buf_splitterG7ton117n243_splitterG7ton242n243_5 , buf_splitterG7ton117n243_splitterG7ton242n243_4 , buf_splitterG7ton117n243_splitterG7ton242n243_3 , buf_splitterG7ton117n243_splitterG7ton242n243_2 , buf_splitterG7ton117n243_splitterG7ton242n243_1 , buf_splitterG8ton159n246_splitterG8ton245n246_10 , buf_splitterG8ton159n246_splitterG8ton245n246_9 , buf_splitterG8ton159n246_splitterG8ton245n246_8 , buf_splitterG8ton159n246_splitterG8ton245n246_7 , buf_splitterG8ton159n246_splitterG8ton245n246_6 , buf_splitterG8ton159n246_splitterG8ton245n246_5 , buf_splitterG8ton159n246_splitterG8ton245n246_4 , buf_splitterG8ton159n246_splitterG8ton245n246_3 , buf_splitterG8ton159n246_splitterG8ton245n246_2 , buf_splitterG8ton159n246_splitterG8ton245n246_1 , buf_splitterG9ton103n250_splitterG9ton58n250_1 , buf_splitterG9ton58n250_splitterG9ton249n250_10 , buf_splitterG9ton58n250_splitterG9ton249n250_9 , buf_splitterG9ton58n250_splitterG9ton249n250_8 , buf_splitterG9ton58n250_splitterG9ton249n250_7 , buf_splitterG9ton58n250_splitterG9ton249n250_6 , buf_splitterG9ton58n250_splitterG9ton249n250_5 , buf_splitterG9ton58n250_splitterG9ton249n250_4 , buf_splitterG9ton58n250_splitterG9ton249n250_3 , buf_splitterG9ton58n250_splitterG9ton249n250_2 , buf_splitterG9ton58n250_splitterG9ton249n250_1 , buf_splittern35ton78n252_n252_1 , buf_splitterfromn72_n277_8 , buf_splitterfromn72_n277_7 , buf_splitterfromn72_n277_6 , buf_splitterfromn72_n277_5 , buf_splitterfromn72_n277_4 , buf_splitterfromn72_n277_3 , buf_splitterfromn72_n277_2 , buf_splitterfromn72_n277_1 , buf_splittern73ton75n278_n278_6 , buf_splittern73ton75n278_n278_5 , buf_splittern73ton75n278_n278_4 , buf_splittern73ton75n278_n278_3 , buf_splittern73ton75n278_n278_2 , buf_splittern73ton75n278_n278_1 , buf_splittern74ton75n275_n275_6 , buf_splittern74ton75n275_n275_5 , buf_splittern74ton75n275_n275_4 , buf_splittern74ton75n275_n275_3 , buf_splittern74ton75n275_n275_2 , buf_splittern74ton75n275_n275_1 , buf_splittern77ton271n253_n253_1 , buf_splitterfromn98_n321_7 , buf_splitterfromn98_n321_6 , buf_splitterfromn98_n321_5 , buf_splitterfromn98_n321_4 , buf_splitterfromn98_n321_3 , buf_splitterfromn98_n321_2 , buf_splitterfromn98_n321_1 , buf_splittern105ton106n309_splittern105ton308n309_2 , buf_splittern105ton106n309_splittern105ton308n309_1 , buf_splitterfromn125_n297_8 , buf_splitterfromn125_n297_7 , buf_splitterfromn125_n297_6 , buf_splitterfromn125_n297_5 , buf_splitterfromn125_n297_4 , buf_splitterfromn125_n297_3 , buf_splitterfromn125_n297_2 , buf_splitterfromn125_n297_1 , buf_splittern128ton129n295_n295_2 , buf_splittern128ton129n295_n295_1 , buf_splitterfromn151_n289_8 , buf_splitterfromn151_n289_7 , buf_splitterfromn151_n289_6 , buf_splitterfromn151_n289_5 , buf_splitterfromn151_n289_4 , buf_splitterfromn151_n289_3 , buf_splitterfromn151_n289_2 , buf_splitterfromn151_n289_1 , buf_splitterfromn171_n293_8 , buf_splitterfromn171_n293_7 , buf_splitterfromn171_n293_6 , buf_splitterfromn171_n293_5 , buf_splitterfromn171_n293_4 , buf_splitterfromn171_n293_3 , buf_splitterfromn171_n293_2 , buf_splitterfromn171_n293_1 , buf_splittern177ton197n272_n272_1 , buf_splitterfromn191_n283_8 , buf_splitterfromn191_n283_7 , buf_splitterfromn191_n283_6 , buf_splitterfromn191_n283_5 , buf_splitterfromn191_n283_4 , buf_splitterfromn191_n283_3 , buf_splitterfromn191_n283_2 , buf_splitterfromn191_n283_1 , buf_splittern192ton193n284_n284_7 , buf_splittern192ton193n284_n284_6 , buf_splittern192ton193n284_n284_5 , buf_splittern192ton193n284_n284_4 , buf_splittern192ton193n284_n284_3 , buf_splittern192ton193n284_n284_2 , buf_splittern192ton193n284_n284_1 , buf_splitterfromn199_n202_2 , buf_splitterfromn199_n202_1 , buf_splittern203ton204n298_splittern203ton321n298_5 , buf_splittern203ton204n298_splittern203ton321n298_4 , buf_splittern203ton204n298_splittern203ton321n298_3 , buf_splittern203ton204n298_splittern203ton321n298_2 , buf_splittern203ton204n298_splittern203ton321n298_1 , buf_splittern203ton279n298_n279_1 , buf_splitterfromn219_n220_3 , buf_splitterfromn219_n220_2 , buf_splitterfromn219_n220_1 , splitterG1ton48n208 , splitterG1ton49n208 , splitterG1ton207n208 , splitterG10ton61n224 , splitterG10ton120n224 , splitterG10ton223n224 , splitterG11ton134n256 , splitterG11ton135n256 , splitterG11ton255n256 , splitterG12ton163n259 , splitterG12ton164n259 , splitterG12ton258n259 , splitterG13ton79n262 , splitterG13ton111n262 , splitterG13ton261n262 , splitterG14ton180n265 , splitterG14ton103n265 , splitterG14ton264n265 , splitterG15ton134n227 , splitterG15ton135n227 , splitterG15ton226n227 , splitterG16ton64n230 , splitterG16ton65n230 , splitterG16ton229n230 , splitterfromG17 , splitterfromG18 , splitterfromG19 , splitterG2ton45n211 , splitterG2ton146n211 , splitterG2ton210n211 , splitterfromG20 , splitterfromG21 , splitterfromG22 , splitterG23ton109n200 , splitterG23ton127n200 , splitterG24ton88n200 , splitterG24ton34n200 , splitterG25ton193n281 , splitterG26ton100n320 , splitterG27ton153n287 , splitterG28ton173n291 , splitterfromG29 , splitterG3ton45n214 , splitterG3ton156n214 , splitterG3ton213n214 , splitterfromG30 , splitterG31ton127n282 , splitterG31ton126n282 , splitterG31ton172n282 , splitterG31ton201n282 , splitterG31ton287n282 , splitterG31ton291n282 , splitterG31ton276n282 , splitterfromG32 , splitterG33ton109n316 , splitterG33ton179n316 , splitterG33ton199n316 , splitterG33ton203n316 , splitterG33ton273n316 , splitterG4ton180n217 , splitterG4ton181n217 , splitterG4ton118n217 , splitterG4ton216n217 , splitterG5ton143n237 , splitterG5ton39n237 , splitterG5ton236n237 , splitterG6ton36n240 , splitterG6ton156n240 , splitterG6ton239n240 , splitterG7ton36n243 , splitterG7ton117n243 , splitterG7ton242n243 , splitterG8ton143n246 , splitterG8ton144n246 , splitterG8ton159n246 , splitterG8ton245n246 , splitterG9ton103n250 , splitterG9ton58n250 , splitterG9ton249n250 , splitterfromn34 , splittern35ton269n252 , splittern35ton78n252 , splitterfromn38 , splittern41ton93n55 , splittern41ton54n55 , splitterfromn44 , splitterfromn47 , splittern50ton51n187 , splitterfromn53 , splittern56ton70n299 , splitterfromn57 , splitterfromn60 , splittern63ton163n65 , splittern66ton85n68 , splitterfromn69 , splitterfromn72 , splittern73ton75n278 , splittern74ton75n275 , splittern77ton271n253 , splitterfromn78 , splitterfromn81 , splitterfromn84 , splittern87ton189n97 , splittern87ton308n97 , splitterfromn88 , splitterfromn89 , splitterfromn92 , splitterfromn95 , splitterfromn98 , splitterfromn99 , splittern105ton106n309 , splittern105ton308n309 , splittern108ton114n141 , splitterfromn109 , splitterfromn110 , splitterfromn113 , splitterfromn116 , splitterfromn119 , splitterfromn122 , splitterfromn125 , splitterfromn126 , splitterfromn127 , splittern128ton129n295 , splitterfromn133 , splitterfromn136 , splitterfromn139 , splitterfromn142 , splitterfromn145 , splitterfromn148 , splitterfromn151 , splitterfromn152 , splitterfromn158 , splitterfromn161 , splitterfromn162 , splitterfromn165 , splitterfromn168 , splitterfromn171 , splitterfromn172 , splittern177ton197n272 , splittern178ton269n232 , splittern178ton196n232 , splitterfromn179 , splitterfromn182 , splitterfromn185 , splitterfromn188 , splitterfromn191 , splittern192ton193n284 , splittern195ton196n270 , splitterfromn197 , splitterfromn198 , splitterfromn199 , splitterfromn200 , splitterfromn201 , splittern203ton204n298 , splittern203ton321n298 , splittern203ton279n298 , splittern203ton285n298 , splitterfromn204 , splitterfromn205 , splittern206ton267n217 , splittern206ton207n217 , splittern206ton207n211 , splittern206ton213n217 , splitterfromn219 , splittern221ton222n254 , splittern222ton267n230 , splittern222ton223n230 , splittern222ton226n230 , splitterfromn234 , splittern235ton236n246 , splittern235ton239n240 , splittern235ton242n246 , splitterfromn248 , splittern254ton255n265 , splittern254ton255n259 , splittern254ton261n265 , splittern267ton275n320 , splittern267ton268n320 , splitterfromn275 , splitterfromn281 , splitterfromn299 , splitterfromn300 , splitterfromn304 , splitterfromn311 , splitterfromn312 , splitterfromn316 ;

PI_AQFP G1_( clk_1 , G1 );
PI_AQFP G10_( clk_1 , G10 );
PI_AQFP G11_( clk_1 , G11 );
PI_AQFP G12_( clk_1 , G12 );
PI_AQFP G13_( clk_1 , G13 );
PI_AQFP G14_( clk_1 , G14 );
PI_AQFP G15_( clk_1 , G15 );
PI_AQFP G16_( clk_1 , G16 );
PI_AQFP G17_( clk_1 , G17 );
PI_AQFP G18_( clk_1 , G18 );
PI_AQFP G19_( clk_1 , G19 );
PI_AQFP G2_( clk_1 , G2 );
PI_AQFP G20_( clk_1 , G20 );
PI_AQFP G21_( clk_1 , G21 );
PI_AQFP G22_( clk_1 , G22 );
PI_AQFP G23_( clk_1 , G23 );
PI_AQFP G24_( clk_1 , G24 );
PI_AQFP G25_( clk_1 , G25 );
PI_AQFP G26_( clk_1 , G26 );
PI_AQFP G27_( clk_1 , G27 );
PI_AQFP G28_( clk_1 , G28 );
PI_AQFP G29_( clk_1 , G29 );
PI_AQFP G3_( clk_1 , G3 );
PI_AQFP G30_( clk_1 , G30 );
PI_AQFP G31_( clk_1 , G31 );
PI_AQFP G32_( clk_1 , G32 );
PI_AQFP G33_( clk_1 , G33 );
PI_AQFP G4_( clk_1 , G4 );
PI_AQFP G5_( clk_1 , G5 );
PI_AQFP G6_( clk_1 , G6 );
PI_AQFP G7_( clk_1 , G7 );
PI_AQFP G8_( clk_1 , G8 );
PI_AQFP G9_( clk_1 , G9 );
or_AQFP n34_( clk_6 , splitterG24ton34n200 , splitterG31ton127n282 , 0 , 0 , n34 );
and_AQFP n35_( clk_8 , buf_splitterfromG18_n35_1 , splitterfromn34 , 0 , 0 , n35 );
or_AQFP n36_( clk_4 , splitterG6ton36n240 , splitterG7ton36n243 , 0 , 0 , n36 );
and_AQFP n37_( clk_4 , splitterG6ton36n240 , splitterG7ton36n243 , 0 , 0 , n37 );
and_AQFP n38_( clk_5 , n36 , n37 , 0 , 1 , n38 );
and_AQFP n39_( clk_7 , splitterG5ton39n237 , splitterfromn38 , 0 , 0 , n39 );
or_AQFP n40_( clk_7 , splitterG5ton39n237 , splitterfromn38 , 0 , 0 , n40 );
and_AQFP n41_( clk_8 , n39 , n40 , 1 , 0 , n41 );
or_AQFP n42_( clk_7 , splitterG4ton118n217 , splitterG8ton144n246 , 0 , 0 , n42 );
and_AQFP n43_( clk_7 , splitterG4ton118n217 , splitterG8ton144n246 , 0 , 0 , n43 );
and_AQFP n44_( clk_8 , n42 , n43 , 0 , 1 , n44 );
or_AQFP n45_( clk_4 , splitterG2ton45n211 , splitterG3ton45n214 , 0 , 0 , n45 );
and_AQFP n46_( clk_4 , splitterG2ton45n211 , splitterG3ton45n214 , 0 , 0 , n46 );
and_AQFP n47_( clk_5 , n45 , n46 , 0 , 1 , n47 );
and_AQFP n48_( clk_7 , buf_splitterG1ton48n208_n48_1 , splitterfromn47 , 0 , 0 , n48 );
or_AQFP n49_( clk_7 , splitterG1ton49n208 , splitterfromn47 , 0 , 0 , n49 );
and_AQFP n50_( clk_8 , n48 , n49 , 1 , 0 , n50 );
and_AQFP n51_( clk_2 , splitterfromn44 , splittern50ton51n187 , 1 , 0 , n51 );
and_AQFP n52_( clk_2 , splitterfromn44 , splittern50ton51n187 , 0 , 1 , n52 );
or_AQFP n53_( clk_3 , n51 , n52 , 0 , 0 , n53 );
or_AQFP n54_( clk_5 , splittern41ton54n55 , splitterfromn53 , 0 , 0 , n54 );
and_AQFP n55_( clk_5 , splittern41ton54n55 , splitterfromn53 , 0 , 0 , n55 );
and_AQFP n56_( clk_6 , n54 , n55 , 0 , 1 , n56 );
and_AQFP n57_( clk_6 , splitterfromG21 , splitterG33ton179n316 , 0 , 1 , n57 );
and_AQFP n58_( clk_8 , splitterG9ton58n250 , splitterfromn57 , 1 , 0 , n58 );
and_AQFP n59_( clk_8 , splitterG9ton58n250 , splitterfromn57 , 0 , 1 , n59 );
or_AQFP n60_( clk_1 , n58 , n59 , 0 , 0 , n60 );
and_AQFP n61_( clk_4 , splitterG10ton61n224 , splitterG15ton135n227 , 0 , 1 , n61 );
and_AQFP n62_( clk_4 , splitterG10ton61n224 , splitterG15ton135n227 , 1 , 0 , n62 );
or_AQFP n63_( clk_5 , n61 , n62 , 0 , 0 , n63 );
and_AQFP n64_( clk_7 , buf_splitterG16ton64n230_n64_1 , splittern63ton163n65 , 1 , 0 , n64 );
and_AQFP n65_( clk_7 , splitterG16ton65n230 , splittern63ton163n65 , 0 , 1 , n65 );
or_AQFP n66_( clk_8 , n64 , n65 , 0 , 0 , n66 );
and_AQFP n67_( clk_3 , splitterfromn60 , splittern66ton85n68 , 1 , 0 , n67 );
and_AQFP n68_( clk_3 , splitterfromn60 , splittern66ton85n68 , 0 , 1 , n68 );
or_AQFP n69_( clk_4 , n67 , n68 , 0 , 0 , n69 );
and_AQFP n70_( clk_8 , splittern56ton70n299 , splitterfromn69 , 0 , 1 , n70 );
and_AQFP n71_( clk_8 , splittern56ton70n299 , splitterfromn69 , 1 , 0 , n71 );
or_AQFP n72_( clk_1 , n70 , n71 , 0 , 0 , n72 );
or_AQFP n73_( clk_3 , splitterG31ton201n282 , splitterfromn72 , 0 , 0 , n73 );
and_AQFP n74_( clk_8 , buf_splitterfromG17_n74_1 , splitterfromn34 , 0 , 0 , n74 );
and_AQFP n75_( clk_5 , splittern73ton75n278 , splittern74ton75n275 , 0 , 1 , n75 );
and_AQFP n76_( clk_5 , splittern73ton75n278 , splittern74ton75n275 , 1 , 0 , n76 );
or_AQFP n77_( clk_6 , n75 , n76 , 0 , 0 , n77 );
and_AQFP n78_( clk_8 , splittern35ton78n252 , splittern77ton271n253 , 0 , 1 , n78 );
and_AQFP n79_( clk_4 , splitterG11ton135n256 , splitterG13ton79n262 , 1 , 0 , n79 );
and_AQFP n80_( clk_4 , splitterG11ton135n256 , splitterG13ton79n262 , 0 , 1 , n80 );
or_AQFP n81_( clk_5 , n79 , n80 , 0 , 0 , n81 );
and_AQFP n82_( clk_7 , splitterG12ton164n259 , splitterfromn81 , 0 , 1 , n82 );
and_AQFP n83_( clk_7 , splitterG12ton164n259 , splitterfromn81 , 1 , 0 , n83 );
or_AQFP n84_( clk_8 , n82 , n83 , 0 , 0 , n84 );
and_AQFP n85_( clk_2 , splittern66ton85n68 , splitterfromn84 , 1 , 0 , n85 );
and_AQFP n86_( clk_2 , splittern66ton85n68 , splitterfromn84 , 0 , 1 , n86 );
or_AQFP n87_( clk_3 , n85 , n86 , 0 , 0 , n87 );
or_AQFP n88_( clk_4 , splitterG24ton88n200 , splitterG33ton109n316 , 0 , 0 , n88 );
and_AQFP n89_( clk_6 , splitterfromG17 , splitterfromn88 , 0 , 1 , n89 );
and_AQFP n90_( clk_8 , splitterG1ton49n208 , splitterfromn89 , 1 , 0 , n90 );
and_AQFP n91_( clk_8 , splitterG1ton49n208 , splitterfromn89 , 0 , 1 , n91 );
or_AQFP n92_( clk_1 , n90 , n91 , 0 , 0 , n92 );
or_AQFP n93_( clk_3 , splittern41ton93n55 , splitterfromn92 , 0 , 0 , n93 );
and_AQFP n94_( clk_3 , splittern41ton93n55 , splitterfromn92 , 0 , 0 , n94 );
and_AQFP n95_( clk_4 , n93 , n94 , 0 , 1 , n95 );
or_AQFP n96_( clk_6 , splittern87ton308n97 , splitterfromn95 , 0 , 0 , n96 );
and_AQFP n97_( clk_6 , splittern87ton308n97 , splitterfromn95 , 0 , 0 , n97 );
and_AQFP n98_( clk_7 , n96 , n97 , 0 , 1 , n98 );
or_AQFP n99_( clk_1 , splitterG31ton172n282 , splitterfromn98 , 0 , 0 , n99 );
or_AQFP n100_( clk_3 , splitterG26ton100n320 , splitterfromn99 , 0 , 0 , n100 );
and_AQFP n101_( clk_3 , splitterG26ton100n320 , splitterfromn99 , 0 , 0 , n101 );
and_AQFP n102_( clk_4 , n100 , n101 , 0 , 1 , n102 );
and_AQFP n103_( clk_5 , splitterG14ton103n265 , splitterG9ton103n250 , 1 , 0 , n103 );
and_AQFP n104_( clk_5 , splitterG14ton103n265 , splitterG9ton103n250 , 0 , 1 , n104 );
or_AQFP n105_( clk_6 , n103 , n104 , 0 , 0 , n105 );
and_AQFP n106_( clk_8 , splitterG16ton65n230 , splittern105ton106n309 , 1 , 0 , n106 );
and_AQFP n107_( clk_8 , splitterG16ton65n230 , splittern105ton106n309 , 0 , 1 , n107 );
or_AQFP n108_( clk_1 , n106 , n107 , 0 , 0 , n108 );
or_AQFP n109_( clk_4 , splitterG23ton109n200 , splitterG33ton109n316 , 0 , 0 , n109 );
and_AQFP n110_( clk_6 , splitterfromG20 , splitterfromn109 , 0 , 1 , n110 );
and_AQFP n111_( clk_8 , splitterG13ton111n262 , splitterfromn110 , 1 , 0 , n111 );
and_AQFP n112_( clk_8 , splitterG13ton111n262 , splitterfromn110 , 0 , 1 , n112 );
or_AQFP n113_( clk_1 , n111 , n112 , 0 , 0 , n113 );
and_AQFP n114_( clk_3 , splittern108ton114n141 , splitterfromn113 , 1 , 0 , n114 );
and_AQFP n115_( clk_3 , splittern108ton114n141 , splitterfromn113 , 0 , 1 , n115 );
or_AQFP n116_( clk_4 , n114 , n115 , 0 , 0 , n116 );
and_AQFP n117_( clk_6 , splitterG4ton181n217 , splitterG7ton117n243 , 0 , 1 , n117 );
and_AQFP n118_( clk_7 , splitterG4ton118n217 , splitterG7ton117n243 , 1 , 0 , n118 );
or_AQFP n119_( clk_8 , n117 , n118 , 0 , 0 , n119 );
and_AQFP n120_( clk_2 , splitterG10ton120n224 , splitterfromn119 , 0 , 1 , n120 );
and_AQFP n121_( clk_2 , splitterG10ton120n224 , splitterfromn119 , 1 , 0 , n121 );
or_AQFP n122_( clk_3 , n120 , n121 , 0 , 0 , n122 );
and_AQFP n123_( clk_6 , splitterfromn116 , splitterfromn122 , 0 , 0 , n123 );
or_AQFP n124_( clk_6 , splitterfromn116 , splitterfromn122 , 0 , 0 , n124 );
and_AQFP n125_( clk_7 , n123 , n124 , 1 , 0 , n125 );
or_AQFP n126_( clk_1 , splitterG31ton126n282 , splitterfromn125 , 0 , 0 , n126 );
or_AQFP n127_( clk_6 , splitterG23ton127n200 , splitterG31ton127n282 , 0 , 0 , n127 );
and_AQFP n128_( clk_8 , buf_splitterfromG19_n128_1 , splitterfromn127 , 0 , 0 , n128 );
and_AQFP n129_( clk_3 , splitterfromn126 , splittern128ton129n295 , 0 , 0 , n129 );
or_AQFP n130_( clk_3 , splitterfromn126 , splittern128ton129n295 , 0 , 0 , n130 );
and_AQFP n131_( clk_4 , n129 , n130 , 1 , 0 , n131 );
and_AQFP n132_( clk_5 , n102 , n131 , 0 , 0 , n132 );
and_AQFP n133_( clk_6 , splitterfromG18 , splitterfromn88 , 0 , 1 , n133 );
or_AQFP n134_( clk_3 , splitterG11ton134n256 , splitterG15ton134n227 , 0 , 0 , n134 );
and_AQFP n135_( clk_4 , splitterG11ton135n256 , splitterG15ton135n227 , 0 , 0 , n135 );
and_AQFP n136_( clk_5 , n134 , n135 , 0 , 1 , n136 );
or_AQFP n137_( clk_8 , splitterfromn133 , splitterfromn136 , 0 , 0 , n137 );
and_AQFP n138_( clk_8 , splitterfromn133 , splitterfromn136 , 0 , 0 , n138 );
and_AQFP n139_( clk_1 , n137 , n138 , 0 , 1 , n139 );
and_AQFP n140_( clk_3 , splittern108ton114n141 , splitterfromn139 , 0 , 0 , n140 );
or_AQFP n141_( clk_3 , splittern108ton114n141 , splitterfromn139 , 0 , 0 , n141 );
and_AQFP n142_( clk_4 , n140 , n141 , 1 , 0 , n142 );
and_AQFP n143_( clk_5 , splitterG5ton143n237 , splitterG8ton143n246 , 0 , 1 , n143 );
and_AQFP n144_( clk_6 , splitterG5ton143n237 , splitterG8ton144n246 , 1 , 0 , n144 );
or_AQFP n145_( clk_7 , n143 , n144 , 0 , 0 , n145 );
and_AQFP n146_( clk_1 , splitterG2ton146n211 , splitterfromn145 , 0 , 1 , n146 );
and_AQFP n147_( clk_1 , splitterG2ton146n211 , splitterfromn145 , 1 , 0 , n147 );
or_AQFP n148_( clk_2 , n146 , n147 , 0 , 0 , n148 );
and_AQFP n149_( clk_6 , splitterfromn142 , splitterfromn148 , 1 , 0 , n149 );
and_AQFP n150_( clk_6 , splitterfromn142 , splitterfromn148 , 0 , 1 , n150 );
or_AQFP n151_( clk_7 , n149 , n150 , 0 , 0 , n151 );
and_AQFP n152_( clk_1 , splitterG31ton126n282 , splitterfromn151 , 1 , 0 , n152 );
and_AQFP n153_( clk_3 , splitterG27ton153n287 , splitterfromn152 , 0 , 0 , n153 );
or_AQFP n154_( clk_3 , splitterG27ton153n287 , splitterfromn152 , 0 , 0 , n154 );
and_AQFP n155_( clk_4 , n153 , n154 , 1 , 0 , n155 );
or_AQFP n156_( clk_6 , splitterG3ton156n214 , splitterG6ton156n240 , 0 , 0 , n156 );
and_AQFP n157_( clk_6 , splitterG3ton156n214 , splitterG6ton156n240 , 0 , 0 , n157 );
and_AQFP n158_( clk_7 , n156 , n157 , 0 , 1 , n158 );
and_AQFP n159_( clk_1 , splitterG8ton159n246 , splitterfromn158 , 0 , 0 , n159 );
or_AQFP n160_( clk_1 , splitterG8ton159n246 , splitterfromn158 , 0 , 0 , n160 );
and_AQFP n161_( clk_2 , n159 , n160 , 1 , 0 , n161 );
and_AQFP n162_( clk_6 , splitterfromG19 , splitterfromn109 , 0 , 1 , n162 );
and_AQFP n163_( clk_7 , buf_splitterG12ton163n259_n163_1 , splittern63ton163n65 , 0 , 0 , n163 );
or_AQFP n164_( clk_7 , splitterG12ton164n259 , splittern63ton163n65 , 0 , 0 , n164 );
and_AQFP n165_( clk_8 , n163 , n164 , 1 , 0 , n165 );
and_AQFP n166_( clk_2 , splitterfromn162 , splitterfromn165 , 0 , 1 , n166 );
and_AQFP n167_( clk_2 , splitterfromn162 , splitterfromn165 , 1 , 0 , n167 );
or_AQFP n168_( clk_3 , n166 , n167 , 0 , 0 , n168 );
or_AQFP n169_( clk_5 , splitterfromn161 , splitterfromn168 , 0 , 0 , n169 );
and_AQFP n170_( clk_5 , splitterfromn161 , splitterfromn168 , 0 , 0 , n170 );
and_AQFP n171_( clk_6 , n169 , n170 , 0 , 1 , n171 );
and_AQFP n172_( clk_1 , splitterG31ton172n282 , splitterfromn171 , 1 , 0 , n172 );
and_AQFP n173_( clk_3 , splitterG28ton173n291 , splitterfromn172 , 0 , 0 , n173 );
or_AQFP n174_( clk_3 , splitterG28ton173n291 , splitterfromn172 , 0 , 0 , n174 );
and_AQFP n175_( clk_4 , n173 , n174 , 1 , 0 , n175 );
or_AQFP n176_( clk_5 , n155 , n175 , 0 , 0 , n176 );
and_AQFP n177_( clk_6 , n132 , n176 , 0 , 1 , n177 );
and_AQFP n178_( clk_8 , buf_splitterfromG20_n178_1 , splitterfromn127 , 0 , 0 , n178 );
and_AQFP n179_( clk_6 , splitterfromG22 , splitterG33ton179n316 , 0 , 1 , n179 );
and_AQFP n180_( clk_4 , splitterG14ton180n265 , splitterG4ton180n217 , 1 , 0 , n180 );
and_AQFP n181_( clk_5 , splitterG14ton103n265 , splitterG4ton181n217 , 0 , 1 , n181 );
or_AQFP n182_( clk_6 , n180 , n181 , 0 , 0 , n182 );
and_AQFP n183_( clk_8 , splitterfromn179 , splitterfromn182 , 0 , 1 , n183 );
and_AQFP n184_( clk_8 , splitterfromn179 , splitterfromn182 , 1 , 0 , n184 );
or_AQFP n185_( clk_1 , n183 , n184 , 0 , 0 , n185 );
or_AQFP n186_( clk_3 , splittern50ton51n187 , splitterfromn185 , 0 , 0 , n186 );
and_AQFP n187_( clk_3 , splittern50ton51n187 , splitterfromn185 , 0 , 0 , n187 );
and_AQFP n188_( clk_4 , n186 , n187 , 0 , 1 , n188 );
or_AQFP n189_( clk_6 , splittern87ton189n97 , splitterfromn188 , 0 , 0 , n189 );
and_AQFP n190_( clk_6 , splittern87ton189n97 , splitterfromn188 , 0 , 0 , n190 );
and_AQFP n191_( clk_7 , n189 , n190 , 0 , 1 , n191 );
and_AQFP n192_( clk_2 , splitterG31ton172n282 , splitterfromn191 , 1 , 0 , n192 );
or_AQFP n193_( clk_4 , splitterG25ton193n281 , splittern192ton193n284 , 0 , 0 , n193 );
and_AQFP n194_( clk_4 , splitterG25ton193n281 , splittern192ton193n284 , 0 , 0 , n194 );
and_AQFP n195_( clk_5 , n193 , n194 , 0 , 1 , n195 );
and_AQFP n196_( clk_7 , splittern178ton196n232 , splittern195ton196n270 , 0 , 0 , n196 );
and_AQFP n197_( clk_8 , splittern177ton197n272 , n196 , 0 , 1 , n197 );
and_AQFP n198_( clk_2 , splitterfromn78 , splitterfromn197 , 1 , 0 , n198 );
or_AQFP n199_( clk_8 , buf_splitterfromG29_n199_1 , splitterG33ton199n316 , 0 , 0 , n199 );
and_AQFP n200_( clk_7 , splitterG23ton127n200 , splitterG24ton34n200 , 1 , 0 , n200 );
or_AQFP n201_( clk_3 , splitterG31ton201n282 , splitterfromn200 , 0 , 0 , n201 );
or_AQFP n202_( clk_5 , buf_splitterfromn199_n202_1 , splitterfromn201 , 0 , 0 , n202 );
or_AQFP n203_( clk_8 , splitterfromG32 , splitterG33ton203n316 , 0 , 0 , n203 );
or_AQFP n204_( clk_3 , splitterfromn200 , splittern203ton204n298 , 0 , 0 , n204 );
and_AQFP n205_( clk_7 , n202 , splitterfromn204 , 0 , 0 , n205 );
and_AQFP n206_( clk_4 , splitterfromn198 , splitterfromn205 , 0 , 1 , n206 );
or_AQFP n207_( clk_8 , splitterG1ton207n208 , splittern206ton207n211 , 0 , 0 , n207 );
and_AQFP n208_( clk_8 , splitterG1ton207n208 , splittern206ton207n211 , 0 , 0 , n208 );
and_AQFP n209_( clk_2 , n207 , n208 , 0 , 1 , n209 );
or_AQFP n210_( clk_8 , splitterG2ton210n211 , splittern206ton207n211 , 0 , 0 , n210 );
and_AQFP n211_( clk_8 , splitterG2ton210n211 , splittern206ton207n211 , 0 , 0 , n211 );
and_AQFP n212_( clk_2 , n210 , n211 , 0 , 1 , n212 );
or_AQFP n213_( clk_8 , splitterG3ton213n214 , splittern206ton213n217 , 0 , 0 , n213 );
and_AQFP n214_( clk_8 , splitterG3ton213n214 , splittern206ton213n217 , 0 , 0 , n214 );
and_AQFP n215_( clk_2 , n213 , n214 , 0 , 1 , n215 );
or_AQFP n216_( clk_8 , splitterG4ton216n217 , splittern206ton213n217 , 0 , 0 , n216 );
and_AQFP n217_( clk_8 , splitterG4ton216n217 , splittern206ton213n217 , 0 , 0 , n217 );
and_AQFP n218_( clk_2 , n216 , n217 , 0 , 1 , n218 );
or_AQFP n219_( clk_8 , buf_splitterfromG30_n219_1 , splitterG33ton199n316 , 0 , 0 , n219 );
or_AQFP n220_( clk_5 , splitterfromn201 , buf_splitterfromn219_n220_1 , 0 , 0 , n220 );
and_AQFP n221_( clk_7 , splitterfromn204 , n220 , 0 , 0 , n221 );
and_AQFP n222_( clk_4 , splitterfromn198 , splittern221ton222n254 , 0 , 1 , n222 );
or_AQFP n223_( clk_7 , splitterG10ton223n224 , splittern222ton223n230 , 0 , 0 , n223 );
and_AQFP n224_( clk_7 , splitterG10ton223n224 , splittern222ton223n230 , 0 , 0 , n224 );
and_AQFP n225_( clk_1 , n223 , n224 , 0 , 1 , n225 );
or_AQFP n226_( clk_8 , splitterG15ton226n227 , splittern222ton226n230 , 0 , 0 , n226 );
and_AQFP n227_( clk_8 , splitterG15ton226n227 , splittern222ton226n230 , 0 , 0 , n227 );
and_AQFP n228_( clk_2 , n226 , n227 , 0 , 1 , n228 );
or_AQFP n229_( clk_8 , splitterG16ton229n230 , splittern222ton226n230 , 0 , 0 , n229 );
and_AQFP n230_( clk_8 , splitterG16ton229n230 , splittern222ton226n230 , 0 , 0 , n230 );
and_AQFP n231_( clk_2 , n229 , n230 , 0 , 1 , n231 );
and_AQFP n232_( clk_7 , splittern178ton196n232 , splittern195ton196n270 , 0 , 1 , n232 );
and_AQFP n233_( clk_8 , splittern177ton197n272 , n232 , 0 , 0 , n233 );
and_AQFP n234_( clk_2 , splitterfromn78 , n233 , 1 , 0 , n234 );
and_AQFP n235_( clk_4 , splitterfromn205 , splitterfromn234 , 1 , 0 , n235 );
or_AQFP n236_( clk_6 , splitterG5ton236n237 , splittern235ton236n246 , 0 , 0 , n236 );
and_AQFP n237_( clk_6 , splitterG5ton236n237 , splittern235ton236n246 , 0 , 0 , n237 );
and_AQFP n238_( clk_8 , n236 , n237 , 0 , 1 , n238 );
or_AQFP n239_( clk_7 , splitterG6ton239n240 , splittern235ton239n240 , 0 , 0 , n239 );
and_AQFP n240_( clk_7 , splitterG6ton239n240 , splittern235ton239n240 , 0 , 0 , n240 );
and_AQFP n241_( clk_1 , n239 , n240 , 0 , 1 , n241 );
or_AQFP n242_( clk_7 , splitterG7ton242n243 , splittern235ton242n246 , 0 , 0 , n242 );
and_AQFP n243_( clk_7 , splitterG7ton242n243 , splittern235ton242n246 , 0 , 0 , n243 );
and_AQFP n244_( clk_1 , n242 , n243 , 0 , 1 , n244 );
or_AQFP n245_( clk_7 , splitterG8ton245n246 , splittern235ton242n246 , 0 , 0 , n245 );
and_AQFP n246_( clk_7 , splitterG8ton245n246 , splittern235ton242n246 , 0 , 0 , n246 );
and_AQFP n247_( clk_1 , n245 , n246 , 0 , 1 , n247 );
and_AQFP n248_( clk_4 , splittern221ton222n254 , splitterfromn234 , 1 , 0 , n248 );
and_AQFP n249_( clk_6 , splitterG9ton249n250 , splitterfromn248 , 0 , 1 , n249 );
and_AQFP n250_( clk_6 , splitterG9ton249n250 , splitterfromn248 , 1 , 0 , n250 );
or_AQFP n251_( clk_8 , n249 , n250 , 0 , 0 , n251 );
and_AQFP n252_( clk_2 , buf_splittern35ton78n252_n252_1 , splitterfromn197 , 0 , 0 , n252 );
and_AQFP n253_( clk_3 , buf_splittern77ton271n253_n253_1 , n252 , 0 , 0 , n253 );
and_AQFP n254_( clk_4 , splittern221ton222n254 , n253 , 1 , 0 , n254 );
or_AQFP n255_( clk_7 , splitterG11ton255n256 , splittern254ton255n259 , 0 , 0 , n255 );
and_AQFP n256_( clk_7 , splitterG11ton255n256 , splittern254ton255n259 , 0 , 0 , n256 );
and_AQFP n257_( clk_1 , n255 , n256 , 0 , 1 , n257 );
or_AQFP n258_( clk_7 , splitterG12ton258n259 , splittern254ton255n259 , 0 , 0 , n258 );
and_AQFP n259_( clk_7 , splitterG12ton258n259 , splittern254ton255n259 , 0 , 0 , n259 );
and_AQFP n260_( clk_1 , n258 , n259 , 0 , 1 , n260 );
or_AQFP n261_( clk_7 , splitterG13ton261n262 , splittern254ton261n265 , 0 , 0 , n261 );
and_AQFP n262_( clk_7 , splitterG13ton261n262 , splittern254ton261n265 , 0 , 0 , n262 );
and_AQFP n263_( clk_1 , n261 , n262 , 0 , 1 , n263 );
or_AQFP n264_( clk_7 , splitterG14ton264n265 , splittern254ton261n265 , 0 , 0 , n264 );
and_AQFP n265_( clk_7 , splitterG14ton264n265 , splittern254ton261n265 , 0 , 0 , n265 );
and_AQFP n266_( clk_1 , n264 , n265 , 0 , 1 , n266 );
or_AQFP n267_( clk_6 , splittern206ton267n217 , splittern222ton267n230 , 0 , 0 , n267 );
and_AQFP n268_( clk_1 , buf_splitterfromG32_n268_1 , splittern267ton268n320 , 0 , 0 , n268 );
or_AQFP n269_( clk_5 , splittern35ton269n252 , splittern178ton269n232 , 0 , 0 , n269 );
or_AQFP n270_( clk_7 , splittern195ton196n270 , n269 , 0 , 0 , n270 );
and_AQFP n271_( clk_8 , splittern77ton271n253 , n270 , 0 , 1 , n271 );
and_AQFP n272_( clk_2 , buf_splittern177ton197n272_n272_1 , n271 , 0 , 0 , n272 );
or_AQFP n273_( clk_8 , splitterG33ton273n316 , buf_n272_n273_1 , 0 , 0 , n273 );
or_AQFP n274_( clk_2 , n268 , n273 , 0 , 0 , n274 );
and_AQFP n275_( clk_8 , buf_splittern74ton75n275_n275_1 , splittern267ton275n320 , 0 , 0 , n275 );
and_AQFP n276_( clk_2 , splitterG31ton276n282 , splitterfromn275 , 1 , 0 , n276 );
and_AQFP n277_( clk_3 , buf_splitterfromn72_n277_1 , n276 , 0 , 1 , n277 );
and_AQFP n278_( clk_2 , buf_splittern73ton75n278_n278_1 , splitterfromn275 , 1 , 0 , n278 );
and_AQFP n279_( clk_3 , buf_splittern203ton279n298_n279_1 , n278 , 0 , 1 , n279 );
and_AQFP n280_( clk_4 , n277 , n279 , 1 , 0 , n280 );
and_AQFP n281_( clk_8 , buf_splitterG25ton193n281_n281_1 , splittern267ton275n320 , 0 , 0 , n281 );
and_AQFP n282_( clk_2 , splitterG31ton276n282 , splitterfromn281 , 1 , 0 , n282 );
or_AQFP n283_( clk_3 , buf_splitterfromn191_n283_1 , n282 , 0 , 0 , n283 );
and_AQFP n284_( clk_2 , buf_splittern192ton193n284_n284_1 , splitterfromn281 , 0 , 0 , n284 );
and_AQFP n285_( clk_3 , splittern203ton285n298 , n284 , 0 , 1 , n285 );
and_AQFP n286_( clk_4 , n283 , n285 , 0 , 0 , n286 );
and_AQFP n287_( clk_5 , buf_splitterG27ton153n287_n287_1 , splitterG31ton287n282 , 0 , 1 , n287 );
and_AQFP n288_( clk_8 , splittern267ton275n320 , buf_n287_n288_1 , 0 , 0 , n288 );
and_AQFP n289_( clk_1 , buf_splitterfromn151_n289_1 , n288 , 0 , 1 , n289 );
and_AQFP n290_( clk_3 , splittern203ton285n298 , n289 , 0 , 1 , n290 );
and_AQFP n291_( clk_7 , buf_splitterG28ton173n291_n291_1 , splitterG31ton291n282 , 0 , 1 , n291 );
and_AQFP n292_( clk_1 , splittern267ton268n320 , buf_n291_n292_1 , 0 , 0 , n292 );
and_AQFP n293_( clk_2 , buf_splitterfromn171_n293_1 , n292 , 0 , 1 , n293 );
and_AQFP n294_( clk_3 , splittern203ton285n298 , n293 , 0 , 1 , n294 );
and_AQFP n295_( clk_7 , splitterG31ton291n282 , buf_splittern128ton129n295_n295_1 , 1 , 0 , n295 );
and_AQFP n296_( clk_1 , splittern267ton268n320 , buf_n295_n296_1 , 0 , 0 , n296 );
or_AQFP n297_( clk_2 , buf_splitterfromn125_n297_1 , n296 , 0 , 0 , n297 );
and_AQFP n298_( clk_3 , splittern203ton285n298 , n297 , 0 , 0 , n298 );
and_AQFP n299_( clk_1 , splittern56ton70n299 , splitterfromn199 , 0 , 0 , n299 );
and_AQFP n300_( clk_6 , splitterfromG21 , splitterfromG29 , 0 , 0 , n300 );
or_AQFP n301_( clk_6 , splittern206ton267n217 , splitterfromn300 , 0 , 0 , n301 );
and_AQFP n302_( clk_6 , splittern206ton267n217 , splitterfromn300 , 0 , 0 , n302 );
and_AQFP n303_( clk_7 , n301 , n302 , 0 , 1 , n303 );
or_AQFP n304_( clk_8 , splitterG33ton273n316 , n303 , 0 , 0 , n304 );
and_AQFP n305_( clk_2 , splitterfromn299 , splitterfromn304 , 0 , 0 , n305 );
or_AQFP n306_( clk_2 , splitterfromn299 , splitterfromn304 , 0 , 0 , n306 );
and_AQFP n307_( clk_3 , n305 , n306 , 1 , 0 , n307 );
or_AQFP n308_( clk_6 , splittern87ton308n97 , splittern105ton308n309 , 0 , 0 , n308 );
and_AQFP n309_( clk_6 , splittern87ton308n97 , splittern105ton308n309 , 0 , 0 , n309 );
and_AQFP n310_( clk_7 , splitterfromn219 , n309 , 0 , 1 , n310 );
and_AQFP n311_( clk_8 , n308 , n310 , 0 , 0 , n311 );
and_AQFP n312_( clk_6 , splitterfromG22 , splitterfromG30 , 0 , 0 , n312 );
or_AQFP n313_( clk_6 , splittern222ton267n230 , splitterfromn312 , 0 , 0 , n313 );
and_AQFP n314_( clk_6 , splittern222ton267n230 , splitterfromn312 , 0 , 0 , n314 );
and_AQFP n315_( clk_7 , n313 , n314 , 0 , 1 , n315 );
or_AQFP n316_( clk_8 , splitterG33ton273n316 , n315 , 0 , 0 , n316 );
and_AQFP n317_( clk_2 , splitterfromn311 , splitterfromn316 , 0 , 1 , n317 );
and_AQFP n318_( clk_2 , splitterfromn311 , splitterfromn316 , 1 , 0 , n318 );
or_AQFP n319_( clk_3 , n317 , n318 , 0 , 0 , n319 );
and_AQFP n320_( clk_1 , buf_splitterG26ton100n320_n320_1 , splittern267ton268n320 , 0 , 0 , n320 );
and_AQFP n321_( clk_7 , buf_splitterfromn98_n321_1 , splittern203ton321n298 , 1 , 0 , n321 );
and_AQFP n322_( clk_2 , n320 , buf_n321_n322_1 , 1 , 0 , n322 );
PO_AQFP G1884_( clk_5 , buf_n209_G1884_1 , 1 , G1884 );
PO_AQFP G1885_( clk_5 , buf_n212_G1885_1 , 1 , G1885 );
PO_AQFP G1886_( clk_5 , buf_n215_G1886_1 , 1 , G1886 );
PO_AQFP G1887_( clk_5 , buf_n218_G1887_1 , 1 , G1887 );
PO_AQFP G1888_( clk_5 , buf_n225_G1888_1 , 1 , G1888 );
PO_AQFP G1889_( clk_5 , buf_n228_G1889_1 , 1 , G1889 );
PO_AQFP G1890_( clk_5 , buf_n231_G1890_1 , 1 , G1890 );
PO_AQFP G1891_( clk_5 , buf_n238_G1891_1 , 1 , G1891 );
PO_AQFP G1892_( clk_5 , buf_n241_G1892_1 , 1 , G1892 );
PO_AQFP G1893_( clk_5 , buf_n244_G1893_1 , 1 , G1893 );
PO_AQFP G1894_( clk_5 , buf_n247_G1894_1 , 1 , G1894 );
PO_AQFP G1895_( clk_5 , buf_n251_G1895_1 , 1 , G1895 );
PO_AQFP G1896_( clk_5 , buf_n257_G1896_1 , 1 , G1896 );
PO_AQFP G1897_( clk_5 , buf_n260_G1897_1 , 1 , G1897 );
PO_AQFP G1898_( clk_5 , buf_n263_G1898_1 , 1 , G1898 );
PO_AQFP G1899_( clk_5 , buf_n266_G1899_1 , 1 , G1899 );
PO_AQFP G1900_( clk_5 , buf_n274_G1900_1 , 0 , G1900 );
PO_AQFP G1901_( clk_5 , n280 , 0 , G1901 );
PO_AQFP G1902_( clk_5 , n286 , 0 , G1902 );
PO_AQFP G1903_( clk_5 , n290 , 0 , G1903 );
PO_AQFP G1904_( clk_5 , n294 , 0 , G1904 );
PO_AQFP G1905_( clk_5 , n298 , 0 , G1905 );
PO_AQFP G1906_( clk_5 , n307 , 1 , G1906 );
PO_AQFP G1907_( clk_5 , n319 , 1 , G1907 );
PO_AQFP G1908_( clk_5 , buf_n322_G1908_1 , 0 , G1908 );
buf_AQFP buf_G1_splitterG1ton48n208_1_( clk_3 , G1 , 0 , buf_G1_splitterG1ton48n208_1 );
buf_AQFP buf_G12_splitterG12ton163n259_1_( clk_3 , G12 , 0 , buf_G12_splitterG12ton163n259_1 );
buf_AQFP buf_G16_splitterG16ton64n230_1_( clk_3 , G16 , 0 , buf_G16_splitterG16ton64n230_1 );
buf_AQFP buf_G17_splitterfromG17_1_( clk_3 , G17 , 0 , buf_G17_splitterfromG17_1 );
buf_AQFP buf_G18_splitterfromG18_1_( clk_3 , G18 , 0 , buf_G18_splitterfromG18_1 );
buf_AQFP buf_G19_splitterfromG19_1_( clk_3 , G19 , 0 , buf_G19_splitterfromG19_1 );
buf_AQFP buf_G20_splitterfromG20_1_( clk_3 , G20 , 0 , buf_G20_splitterfromG20_1 );
buf_AQFP buf_G21_splitterfromG21_1_( clk_3 , G21 , 0 , buf_G21_splitterfromG21_1 );
buf_AQFP buf_G22_splitterfromG22_1_( clk_3 , G22 , 0 , buf_G22_splitterfromG22_1 );
buf_AQFP buf_G25_splitterG25ton193n281_8_( clk_3 , G25 , 0 , buf_G25_splitterG25ton193n281_8 );
buf_AQFP buf_G25_splitterG25ton193n281_7_( clk_5 , buf_G25_splitterG25ton193n281_8 , 0 , buf_G25_splitterG25ton193n281_7 );
buf_AQFP buf_G25_splitterG25ton193n281_6_( clk_7 , buf_G25_splitterG25ton193n281_7 , 0 , buf_G25_splitterG25ton193n281_6 );
buf_AQFP buf_G25_splitterG25ton193n281_5_( clk_1 , buf_G25_splitterG25ton193n281_6 , 0 , buf_G25_splitterG25ton193n281_5 );
buf_AQFP buf_G25_splitterG25ton193n281_4_( clk_3 , buf_G25_splitterG25ton193n281_5 , 0 , buf_G25_splitterG25ton193n281_4 );
buf_AQFP buf_G25_splitterG25ton193n281_3_( clk_5 , buf_G25_splitterG25ton193n281_4 , 0 , buf_G25_splitterG25ton193n281_3 );
buf_AQFP buf_G25_splitterG25ton193n281_2_( clk_7 , buf_G25_splitterG25ton193n281_3 , 0 , buf_G25_splitterG25ton193n281_2 );
buf_AQFP buf_G25_splitterG25ton193n281_1_( clk_1 , buf_G25_splitterG25ton193n281_2 , 0 , buf_G25_splitterG25ton193n281_1 );
buf_AQFP buf_G26_splitterG26ton100n320_7_( clk_3 , G26 , 0 , buf_G26_splitterG26ton100n320_7 );
buf_AQFP buf_G26_splitterG26ton100n320_6_( clk_5 , buf_G26_splitterG26ton100n320_7 , 0 , buf_G26_splitterG26ton100n320_6 );
buf_AQFP buf_G26_splitterG26ton100n320_5_( clk_7 , buf_G26_splitterG26ton100n320_6 , 0 , buf_G26_splitterG26ton100n320_5 );
buf_AQFP buf_G26_splitterG26ton100n320_4_( clk_1 , buf_G26_splitterG26ton100n320_5 , 0 , buf_G26_splitterG26ton100n320_4 );
buf_AQFP buf_G26_splitterG26ton100n320_3_( clk_3 , buf_G26_splitterG26ton100n320_4 , 0 , buf_G26_splitterG26ton100n320_3 );
buf_AQFP buf_G26_splitterG26ton100n320_2_( clk_5 , buf_G26_splitterG26ton100n320_3 , 0 , buf_G26_splitterG26ton100n320_2 );
buf_AQFP buf_G26_splitterG26ton100n320_1_( clk_7 , buf_G26_splitterG26ton100n320_2 , 0 , buf_G26_splitterG26ton100n320_1 );
buf_AQFP buf_G27_splitterG27ton153n287_7_( clk_3 , G27 , 0 , buf_G27_splitterG27ton153n287_7 );
buf_AQFP buf_G27_splitterG27ton153n287_6_( clk_5 , buf_G27_splitterG27ton153n287_7 , 0 , buf_G27_splitterG27ton153n287_6 );
buf_AQFP buf_G27_splitterG27ton153n287_5_( clk_7 , buf_G27_splitterG27ton153n287_6 , 0 , buf_G27_splitterG27ton153n287_5 );
buf_AQFP buf_G27_splitterG27ton153n287_4_( clk_1 , buf_G27_splitterG27ton153n287_5 , 0 , buf_G27_splitterG27ton153n287_4 );
buf_AQFP buf_G27_splitterG27ton153n287_3_( clk_3 , buf_G27_splitterG27ton153n287_4 , 0 , buf_G27_splitterG27ton153n287_3 );
buf_AQFP buf_G27_splitterG27ton153n287_2_( clk_5 , buf_G27_splitterG27ton153n287_3 , 0 , buf_G27_splitterG27ton153n287_2 );
buf_AQFP buf_G27_splitterG27ton153n287_1_( clk_7 , buf_G27_splitterG27ton153n287_2 , 0 , buf_G27_splitterG27ton153n287_1 );
buf_AQFP buf_G28_splitterG28ton173n291_7_( clk_3 , G28 , 0 , buf_G28_splitterG28ton173n291_7 );
buf_AQFP buf_G28_splitterG28ton173n291_6_( clk_5 , buf_G28_splitterG28ton173n291_7 , 0 , buf_G28_splitterG28ton173n291_6 );
buf_AQFP buf_G28_splitterG28ton173n291_5_( clk_7 , buf_G28_splitterG28ton173n291_6 , 0 , buf_G28_splitterG28ton173n291_5 );
buf_AQFP buf_G28_splitterG28ton173n291_4_( clk_1 , buf_G28_splitterG28ton173n291_5 , 0 , buf_G28_splitterG28ton173n291_4 );
buf_AQFP buf_G28_splitterG28ton173n291_3_( clk_3 , buf_G28_splitterG28ton173n291_4 , 0 , buf_G28_splitterG28ton173n291_3 );
buf_AQFP buf_G28_splitterG28ton173n291_2_( clk_5 , buf_G28_splitterG28ton173n291_3 , 0 , buf_G28_splitterG28ton173n291_2 );
buf_AQFP buf_G28_splitterG28ton173n291_1_( clk_7 , buf_G28_splitterG28ton173n291_2 , 0 , buf_G28_splitterG28ton173n291_1 );
buf_AQFP buf_G29_splitterfromG29_1_( clk_3 , G29 , 0 , buf_G29_splitterfromG29_1 );
buf_AQFP buf_G30_splitterfromG30_1_( clk_3 , G30 , 0 , buf_G30_splitterfromG30_1 );
buf_AQFP buf_G31_splitterG31ton127n282_1_( clk_3 , G31 , 0 , buf_G31_splitterG31ton127n282_1 );
buf_AQFP buf_G32_splitterfromG32_6_( clk_3 , G32 , 0 , buf_G32_splitterfromG32_6 );
buf_AQFP buf_G32_splitterfromG32_5_( clk_5 , buf_G32_splitterfromG32_6 , 0 , buf_G32_splitterfromG32_5 );
buf_AQFP buf_G32_splitterfromG32_4_( clk_7 , buf_G32_splitterfromG32_5 , 0 , buf_G32_splitterfromG32_4 );
buf_AQFP buf_G32_splitterfromG32_3_( clk_1 , buf_G32_splitterfromG32_4 , 0 , buf_G32_splitterfromG32_3 );
buf_AQFP buf_G32_splitterfromG32_2_( clk_3 , buf_G32_splitterfromG32_3 , 0 , buf_G32_splitterfromG32_2 );
buf_AQFP buf_G32_splitterfromG32_1_( clk_5 , buf_G32_splitterfromG32_2 , 0 , buf_G32_splitterfromG32_1 );
buf_AQFP buf_G5_splitterG5ton143n237_1_( clk_3 , G5 , 0 , buf_G5_splitterG5ton143n237_1 );
buf_AQFP buf_n35_splittern35ton269n252_5_( clk_2 , n35 , 0 , buf_n35_splittern35ton269n252_5 );
buf_AQFP buf_n35_splittern35ton269n252_4_( clk_4 , buf_n35_splittern35ton269n252_5 , 0 , buf_n35_splittern35ton269n252_4 );
buf_AQFP buf_n35_splittern35ton269n252_3_( clk_6 , buf_n35_splittern35ton269n252_4 , 0 , buf_n35_splittern35ton269n252_3 );
buf_AQFP buf_n35_splittern35ton269n252_2_( clk_8 , buf_n35_splittern35ton269n252_3 , 0 , buf_n35_splittern35ton269n252_2 );
buf_AQFP buf_n35_splittern35ton269n252_1_( clk_2 , buf_n35_splittern35ton269n252_2 , 0 , buf_n35_splittern35ton269n252_1 );
buf_AQFP buf_n74_splittern74ton75n275_5_( clk_2 , n74 , 0 , buf_n74_splittern74ton75n275_5 );
buf_AQFP buf_n74_splittern74ton75n275_4_( clk_4 , buf_n74_splittern74ton75n275_5 , 0 , buf_n74_splittern74ton75n275_4 );
buf_AQFP buf_n74_splittern74ton75n275_3_( clk_6 , buf_n74_splittern74ton75n275_4 , 0 , buf_n74_splittern74ton75n275_3 );
buf_AQFP buf_n74_splittern74ton75n275_2_( clk_8 , buf_n74_splittern74ton75n275_3 , 0 , buf_n74_splittern74ton75n275_2 );
buf_AQFP buf_n74_splittern74ton75n275_1_( clk_2 , buf_n74_splittern74ton75n275_2 , 0 , buf_n74_splittern74ton75n275_1 );
buf_AQFP buf_n128_splittern128ton129n295_4_( clk_2 , n128 , 0 , buf_n128_splittern128ton129n295_4 );
buf_AQFP buf_n128_splittern128ton129n295_3_( clk_4 , buf_n128_splittern128ton129n295_4 , 0 , buf_n128_splittern128ton129n295_3 );
buf_AQFP buf_n128_splittern128ton129n295_2_( clk_6 , buf_n128_splittern128ton129n295_3 , 0 , buf_n128_splittern128ton129n295_2 );
buf_AQFP buf_n128_splittern128ton129n295_1_( clk_8 , buf_n128_splittern128ton129n295_2 , 0 , buf_n128_splittern128ton129n295_1 );
buf_AQFP buf_n178_splittern178ton269n232_5_( clk_2 , n178 , 0 , buf_n178_splittern178ton269n232_5 );
buf_AQFP buf_n178_splittern178ton269n232_4_( clk_4 , buf_n178_splittern178ton269n232_5 , 0 , buf_n178_splittern178ton269n232_4 );
buf_AQFP buf_n178_splittern178ton269n232_3_( clk_6 , buf_n178_splittern178ton269n232_4 , 0 , buf_n178_splittern178ton269n232_3 );
buf_AQFP buf_n178_splittern178ton269n232_2_( clk_8 , buf_n178_splittern178ton269n232_3 , 0 , buf_n178_splittern178ton269n232_2 );
buf_AQFP buf_n178_splittern178ton269n232_1_( clk_2 , buf_n178_splittern178ton269n232_2 , 0 , buf_n178_splittern178ton269n232_1 );
buf_AQFP buf_n199_splitterfromn199_3_( clk_2 , n199 , 0 , buf_n199_splitterfromn199_3 );
buf_AQFP buf_n199_splitterfromn199_2_( clk_4 , buf_n199_splitterfromn199_3 , 0 , buf_n199_splitterfromn199_2 );
buf_AQFP buf_n199_splitterfromn199_1_( clk_6 , buf_n199_splitterfromn199_2 , 0 , buf_n199_splitterfromn199_1 );
buf_AQFP buf_n200_splitterfromn200_4_( clk_1 , n200 , 0 , buf_n200_splitterfromn200_4 );
buf_AQFP buf_n200_splitterfromn200_3_( clk_3 , buf_n200_splitterfromn200_4 , 0 , buf_n200_splitterfromn200_3 );
buf_AQFP buf_n200_splitterfromn200_2_( clk_5 , buf_n200_splitterfromn200_3 , 0 , buf_n200_splitterfromn200_2 );
buf_AQFP buf_n200_splitterfromn200_1_( clk_7 , buf_n200_splitterfromn200_2 , 0 , buf_n200_splitterfromn200_1 );
buf_AQFP buf_n205_splitterfromn205_1_( clk_1 , n205 , 0 , buf_n205_splitterfromn205_1 );
buf_AQFP buf_n209_G1884_1_( clk_4 , n209 , 0 , buf_n209_G1884_1 );
buf_AQFP buf_n212_G1885_1_( clk_4 , n212 , 0 , buf_n212_G1885_1 );
buf_AQFP buf_n215_G1886_1_( clk_4 , n215 , 0 , buf_n215_G1886_1 );
buf_AQFP buf_n218_G1887_1_( clk_4 , n218 , 0 , buf_n218_G1887_1 );
buf_AQFP buf_n219_splitterfromn219_2_( clk_2 , n219 , 0 , buf_n219_splitterfromn219_2 );
buf_AQFP buf_n219_splitterfromn219_1_( clk_4 , buf_n219_splitterfromn219_2 , 0 , buf_n219_splitterfromn219_1 );
buf_AQFP buf_n221_splittern221ton222n254_1_( clk_1 , n221 , 0 , buf_n221_splittern221ton222n254_1 );
buf_AQFP buf_n225_G1888_1_( clk_3 , n225 , 0 , buf_n225_G1888_1 );
buf_AQFP buf_n228_G1889_1_( clk_4 , n228 , 0 , buf_n228_G1889_1 );
buf_AQFP buf_n231_G1890_1_( clk_4 , n231 , 0 , buf_n231_G1890_1 );
buf_AQFP buf_n238_G1891_2_( clk_2 , n238 , 0 , buf_n238_G1891_2 );
buf_AQFP buf_n238_G1891_1_( clk_4 , buf_n238_G1891_2 , 0 , buf_n238_G1891_1 );
buf_AQFP buf_n241_G1892_1_( clk_3 , n241 , 0 , buf_n241_G1892_1 );
buf_AQFP buf_n244_G1893_1_( clk_3 , n244 , 0 , buf_n244_G1893_1 );
buf_AQFP buf_n247_G1894_1_( clk_3 , n247 , 0 , buf_n247_G1894_1 );
buf_AQFP buf_n251_G1895_2_( clk_2 , n251 , 0 , buf_n251_G1895_2 );
buf_AQFP buf_n251_G1895_1_( clk_4 , buf_n251_G1895_2 , 0 , buf_n251_G1895_1 );
buf_AQFP buf_n257_G1896_1_( clk_3 , n257 , 0 , buf_n257_G1896_1 );
buf_AQFP buf_n260_G1897_1_( clk_3 , n260 , 0 , buf_n260_G1897_1 );
buf_AQFP buf_n263_G1898_1_( clk_3 , n263 , 0 , buf_n263_G1898_1 );
buf_AQFP buf_n266_G1899_1_( clk_3 , n266 , 0 , buf_n266_G1899_1 );
buf_AQFP buf_n272_n273_2_( clk_4 , n272 , 0 , buf_n272_n273_2 );
buf_AQFP buf_n272_n273_1_( clk_6 , buf_n272_n273_2 , 0 , buf_n272_n273_1 );
buf_AQFP buf_n274_G1900_1_( clk_4 , n274 , 0 , buf_n274_G1900_1 );
buf_AQFP buf_n287_n288_5_( clk_7 , n287 , 0 , buf_n287_n288_5 );
buf_AQFP buf_n287_n288_4_( clk_1 , buf_n287_n288_5 , 0 , buf_n287_n288_4 );
buf_AQFP buf_n287_n288_3_( clk_3 , buf_n287_n288_4 , 0 , buf_n287_n288_3 );
buf_AQFP buf_n287_n288_2_( clk_5 , buf_n287_n288_3 , 0 , buf_n287_n288_2 );
buf_AQFP buf_n287_n288_1_( clk_7 , buf_n287_n288_2 , 0 , buf_n287_n288_1 );
buf_AQFP buf_n291_n292_4_( clk_1 , n291 , 0 , buf_n291_n292_4 );
buf_AQFP buf_n291_n292_3_( clk_3 , buf_n291_n292_4 , 0 , buf_n291_n292_3 );
buf_AQFP buf_n291_n292_2_( clk_5 , buf_n291_n292_3 , 0 , buf_n291_n292_2 );
buf_AQFP buf_n291_n292_1_( clk_7 , buf_n291_n292_2 , 0 , buf_n291_n292_1 );
buf_AQFP buf_n295_n296_4_( clk_1 , n295 , 0 , buf_n295_n296_4 );
buf_AQFP buf_n295_n296_3_( clk_3 , buf_n295_n296_4 , 0 , buf_n295_n296_3 );
buf_AQFP buf_n295_n296_2_( clk_5 , buf_n295_n296_3 , 0 , buf_n295_n296_2 );
buf_AQFP buf_n295_n296_1_( clk_7 , buf_n295_n296_2 , 0 , buf_n295_n296_1 );
buf_AQFP buf_n299_splitterfromn299_7_( clk_3 , n299 , 0 , buf_n299_splitterfromn299_7 );
buf_AQFP buf_n299_splitterfromn299_6_( clk_5 , buf_n299_splitterfromn299_7 , 0 , buf_n299_splitterfromn299_6 );
buf_AQFP buf_n299_splitterfromn299_5_( clk_7 , buf_n299_splitterfromn299_6 , 0 , buf_n299_splitterfromn299_5 );
buf_AQFP buf_n299_splitterfromn299_4_( clk_1 , buf_n299_splitterfromn299_5 , 0 , buf_n299_splitterfromn299_4 );
buf_AQFP buf_n299_splitterfromn299_3_( clk_3 , buf_n299_splitterfromn299_4 , 0 , buf_n299_splitterfromn299_3 );
buf_AQFP buf_n299_splitterfromn299_2_( clk_5 , buf_n299_splitterfromn299_3 , 0 , buf_n299_splitterfromn299_2 );
buf_AQFP buf_n299_splitterfromn299_1_( clk_7 , buf_n299_splitterfromn299_2 , 0 , buf_n299_splitterfromn299_1 );
buf_AQFP buf_n300_splitterfromn300_10_( clk_8 , n300 , 0 , buf_n300_splitterfromn300_10 );
buf_AQFP buf_n300_splitterfromn300_9_( clk_2 , buf_n300_splitterfromn300_10 , 0 , buf_n300_splitterfromn300_9 );
buf_AQFP buf_n300_splitterfromn300_8_( clk_4 , buf_n300_splitterfromn300_9 , 0 , buf_n300_splitterfromn300_8 );
buf_AQFP buf_n300_splitterfromn300_7_( clk_6 , buf_n300_splitterfromn300_8 , 0 , buf_n300_splitterfromn300_7 );
buf_AQFP buf_n300_splitterfromn300_6_( clk_8 , buf_n300_splitterfromn300_7 , 0 , buf_n300_splitterfromn300_6 );
buf_AQFP buf_n300_splitterfromn300_5_( clk_2 , buf_n300_splitterfromn300_6 , 0 , buf_n300_splitterfromn300_5 );
buf_AQFP buf_n300_splitterfromn300_4_( clk_4 , buf_n300_splitterfromn300_5 , 0 , buf_n300_splitterfromn300_4 );
buf_AQFP buf_n300_splitterfromn300_3_( clk_6 , buf_n300_splitterfromn300_4 , 0 , buf_n300_splitterfromn300_3 );
buf_AQFP buf_n300_splitterfromn300_2_( clk_8 , buf_n300_splitterfromn300_3 , 0 , buf_n300_splitterfromn300_2 );
buf_AQFP buf_n300_splitterfromn300_1_( clk_2 , buf_n300_splitterfromn300_2 , 0 , buf_n300_splitterfromn300_1 );
buf_AQFP buf_n311_splitterfromn311_7_( clk_2 , n311 , 0 , buf_n311_splitterfromn311_7 );
buf_AQFP buf_n311_splitterfromn311_6_( clk_4 , buf_n311_splitterfromn311_7 , 0 , buf_n311_splitterfromn311_6 );
buf_AQFP buf_n311_splitterfromn311_5_( clk_6 , buf_n311_splitterfromn311_6 , 0 , buf_n311_splitterfromn311_5 );
buf_AQFP buf_n311_splitterfromn311_4_( clk_8 , buf_n311_splitterfromn311_5 , 0 , buf_n311_splitterfromn311_4 );
buf_AQFP buf_n311_splitterfromn311_3_( clk_2 , buf_n311_splitterfromn311_4 , 0 , buf_n311_splitterfromn311_3 );
buf_AQFP buf_n311_splitterfromn311_2_( clk_4 , buf_n311_splitterfromn311_3 , 0 , buf_n311_splitterfromn311_2 );
buf_AQFP buf_n311_splitterfromn311_1_( clk_6 , buf_n311_splitterfromn311_2 , 0 , buf_n311_splitterfromn311_1 );
buf_AQFP buf_n312_splitterfromn312_10_( clk_8 , n312 , 0 , buf_n312_splitterfromn312_10 );
buf_AQFP buf_n312_splitterfromn312_9_( clk_2 , buf_n312_splitterfromn312_10 , 0 , buf_n312_splitterfromn312_9 );
buf_AQFP buf_n312_splitterfromn312_8_( clk_4 , buf_n312_splitterfromn312_9 , 0 , buf_n312_splitterfromn312_8 );
buf_AQFP buf_n312_splitterfromn312_7_( clk_6 , buf_n312_splitterfromn312_8 , 0 , buf_n312_splitterfromn312_7 );
buf_AQFP buf_n312_splitterfromn312_6_( clk_8 , buf_n312_splitterfromn312_7 , 0 , buf_n312_splitterfromn312_6 );
buf_AQFP buf_n312_splitterfromn312_5_( clk_2 , buf_n312_splitterfromn312_6 , 0 , buf_n312_splitterfromn312_5 );
buf_AQFP buf_n312_splitterfromn312_4_( clk_4 , buf_n312_splitterfromn312_5 , 0 , buf_n312_splitterfromn312_4 );
buf_AQFP buf_n312_splitterfromn312_3_( clk_6 , buf_n312_splitterfromn312_4 , 0 , buf_n312_splitterfromn312_3 );
buf_AQFP buf_n312_splitterfromn312_2_( clk_8 , buf_n312_splitterfromn312_3 , 0 , buf_n312_splitterfromn312_2 );
buf_AQFP buf_n312_splitterfromn312_1_( clk_2 , buf_n312_splitterfromn312_2 , 0 , buf_n312_splitterfromn312_1 );
buf_AQFP buf_n321_n322_1_( clk_1 , n321 , 0 , buf_n321_n322_1 );
buf_AQFP buf_n322_G1908_1_( clk_4 , n322 , 0 , buf_n322_G1908_1 );
buf_AQFP buf_splitterG1ton48n208_n48_1_( clk_6 , splitterG1ton48n208 , 0 , buf_splitterG1ton48n208_n48_1 );
buf_AQFP buf_splitterG1ton49n208_splitterG1ton207n208_11_( clk_8 , splitterG1ton49n208 , 0 , buf_splitterG1ton49n208_splitterG1ton207n208_11 );
buf_AQFP buf_splitterG1ton49n208_splitterG1ton207n208_10_( clk_2 , buf_splitterG1ton49n208_splitterG1ton207n208_11 , 0 , buf_splitterG1ton49n208_splitterG1ton207n208_10 );
buf_AQFP buf_splitterG1ton49n208_splitterG1ton207n208_9_( clk_4 , buf_splitterG1ton49n208_splitterG1ton207n208_10 , 0 , buf_splitterG1ton49n208_splitterG1ton207n208_9 );
buf_AQFP buf_splitterG1ton49n208_splitterG1ton207n208_8_( clk_6 , buf_splitterG1ton49n208_splitterG1ton207n208_9 , 0 , buf_splitterG1ton49n208_splitterG1ton207n208_8 );
buf_AQFP buf_splitterG1ton49n208_splitterG1ton207n208_7_( clk_8 , buf_splitterG1ton49n208_splitterG1ton207n208_8 , 0 , buf_splitterG1ton49n208_splitterG1ton207n208_7 );
buf_AQFP buf_splitterG1ton49n208_splitterG1ton207n208_6_( clk_2 , buf_splitterG1ton49n208_splitterG1ton207n208_7 , 0 , buf_splitterG1ton49n208_splitterG1ton207n208_6 );
buf_AQFP buf_splitterG1ton49n208_splitterG1ton207n208_5_( clk_4 , buf_splitterG1ton49n208_splitterG1ton207n208_6 , 0 , buf_splitterG1ton49n208_splitterG1ton207n208_5 );
buf_AQFP buf_splitterG1ton49n208_splitterG1ton207n208_4_( clk_6 , buf_splitterG1ton49n208_splitterG1ton207n208_5 , 0 , buf_splitterG1ton49n208_splitterG1ton207n208_4 );
buf_AQFP buf_splitterG1ton49n208_splitterG1ton207n208_3_( clk_8 , buf_splitterG1ton49n208_splitterG1ton207n208_4 , 0 , buf_splitterG1ton49n208_splitterG1ton207n208_3 );
buf_AQFP buf_splitterG1ton49n208_splitterG1ton207n208_2_( clk_2 , buf_splitterG1ton49n208_splitterG1ton207n208_3 , 0 , buf_splitterG1ton49n208_splitterG1ton207n208_2 );
buf_AQFP buf_splitterG1ton49n208_splitterG1ton207n208_1_( clk_4 , buf_splitterG1ton49n208_splitterG1ton207n208_2 , 0 , buf_splitterG1ton49n208_splitterG1ton207n208_1 );
buf_AQFP buf_splitterG10ton61n224_splitterG10ton120n224_2_( clk_5 , splitterG10ton61n224 , 0 , buf_splitterG10ton61n224_splitterG10ton120n224_2 );
buf_AQFP buf_splitterG10ton61n224_splitterG10ton120n224_1_( clk_7 , buf_splitterG10ton61n224_splitterG10ton120n224_2 , 0 , buf_splitterG10ton61n224_splitterG10ton120n224_1 );
buf_AQFP buf_splitterG10ton120n224_splitterG10ton223n224_10_( clk_2 , splitterG10ton120n224 , 0 , buf_splitterG10ton120n224_splitterG10ton223n224_10 );
buf_AQFP buf_splitterG10ton120n224_splitterG10ton223n224_9_( clk_4 , buf_splitterG10ton120n224_splitterG10ton223n224_10 , 0 , buf_splitterG10ton120n224_splitterG10ton223n224_9 );
buf_AQFP buf_splitterG10ton120n224_splitterG10ton223n224_8_( clk_6 , buf_splitterG10ton120n224_splitterG10ton223n224_9 , 0 , buf_splitterG10ton120n224_splitterG10ton223n224_8 );
buf_AQFP buf_splitterG10ton120n224_splitterG10ton223n224_7_( clk_8 , buf_splitterG10ton120n224_splitterG10ton223n224_8 , 0 , buf_splitterG10ton120n224_splitterG10ton223n224_7 );
buf_AQFP buf_splitterG10ton120n224_splitterG10ton223n224_6_( clk_2 , buf_splitterG10ton120n224_splitterG10ton223n224_7 , 0 , buf_splitterG10ton120n224_splitterG10ton223n224_6 );
buf_AQFP buf_splitterG10ton120n224_splitterG10ton223n224_5_( clk_4 , buf_splitterG10ton120n224_splitterG10ton223n224_6 , 0 , buf_splitterG10ton120n224_splitterG10ton223n224_5 );
buf_AQFP buf_splitterG10ton120n224_splitterG10ton223n224_4_( clk_6 , buf_splitterG10ton120n224_splitterG10ton223n224_5 , 0 , buf_splitterG10ton120n224_splitterG10ton223n224_4 );
buf_AQFP buf_splitterG10ton120n224_splitterG10ton223n224_3_( clk_8 , buf_splitterG10ton120n224_splitterG10ton223n224_4 , 0 , buf_splitterG10ton120n224_splitterG10ton223n224_3 );
buf_AQFP buf_splitterG10ton120n224_splitterG10ton223n224_2_( clk_2 , buf_splitterG10ton120n224_splitterG10ton223n224_3 , 0 , buf_splitterG10ton120n224_splitterG10ton223n224_2 );
buf_AQFP buf_splitterG10ton120n224_splitterG10ton223n224_1_( clk_4 , buf_splitterG10ton120n224_splitterG10ton223n224_2 , 0 , buf_splitterG10ton120n224_splitterG10ton223n224_1 );
buf_AQFP buf_splitterG11ton135n256_splitterG11ton255n256_12_( clk_5 , splitterG11ton135n256 , 0 , buf_splitterG11ton135n256_splitterG11ton255n256_12 );
buf_AQFP buf_splitterG11ton135n256_splitterG11ton255n256_11_( clk_7 , buf_splitterG11ton135n256_splitterG11ton255n256_12 , 0 , buf_splitterG11ton135n256_splitterG11ton255n256_11 );
buf_AQFP buf_splitterG11ton135n256_splitterG11ton255n256_10_( clk_1 , buf_splitterG11ton135n256_splitterG11ton255n256_11 , 0 , buf_splitterG11ton135n256_splitterG11ton255n256_10 );
buf_AQFP buf_splitterG11ton135n256_splitterG11ton255n256_9_( clk_3 , buf_splitterG11ton135n256_splitterG11ton255n256_10 , 0 , buf_splitterG11ton135n256_splitterG11ton255n256_9 );
buf_AQFP buf_splitterG11ton135n256_splitterG11ton255n256_8_( clk_5 , buf_splitterG11ton135n256_splitterG11ton255n256_9 , 0 , buf_splitterG11ton135n256_splitterG11ton255n256_8 );
buf_AQFP buf_splitterG11ton135n256_splitterG11ton255n256_7_( clk_7 , buf_splitterG11ton135n256_splitterG11ton255n256_8 , 0 , buf_splitterG11ton135n256_splitterG11ton255n256_7 );
buf_AQFP buf_splitterG11ton135n256_splitterG11ton255n256_6_( clk_1 , buf_splitterG11ton135n256_splitterG11ton255n256_7 , 0 , buf_splitterG11ton135n256_splitterG11ton255n256_6 );
buf_AQFP buf_splitterG11ton135n256_splitterG11ton255n256_5_( clk_3 , buf_splitterG11ton135n256_splitterG11ton255n256_6 , 0 , buf_splitterG11ton135n256_splitterG11ton255n256_5 );
buf_AQFP buf_splitterG11ton135n256_splitterG11ton255n256_4_( clk_5 , buf_splitterG11ton135n256_splitterG11ton255n256_5 , 0 , buf_splitterG11ton135n256_splitterG11ton255n256_4 );
buf_AQFP buf_splitterG11ton135n256_splitterG11ton255n256_3_( clk_7 , buf_splitterG11ton135n256_splitterG11ton255n256_4 , 0 , buf_splitterG11ton135n256_splitterG11ton255n256_3 );
buf_AQFP buf_splitterG11ton135n256_splitterG11ton255n256_2_( clk_1 , buf_splitterG11ton135n256_splitterG11ton255n256_3 , 0 , buf_splitterG11ton135n256_splitterG11ton255n256_2 );
buf_AQFP buf_splitterG11ton135n256_splitterG11ton255n256_1_( clk_3 , buf_splitterG11ton135n256_splitterG11ton255n256_2 , 0 , buf_splitterG11ton135n256_splitterG11ton255n256_1 );
buf_AQFP buf_splitterG12ton163n259_n163_1_( clk_6 , splitterG12ton163n259 , 0 , buf_splitterG12ton163n259_n163_1 );
buf_AQFP buf_splitterG12ton164n259_splitterG12ton258n259_11_( clk_8 , splitterG12ton164n259 , 0 , buf_splitterG12ton164n259_splitterG12ton258n259_11 );
buf_AQFP buf_splitterG12ton164n259_splitterG12ton258n259_10_( clk_2 , buf_splitterG12ton164n259_splitterG12ton258n259_11 , 0 , buf_splitterG12ton164n259_splitterG12ton258n259_10 );
buf_AQFP buf_splitterG12ton164n259_splitterG12ton258n259_9_( clk_4 , buf_splitterG12ton164n259_splitterG12ton258n259_10 , 0 , buf_splitterG12ton164n259_splitterG12ton258n259_9 );
buf_AQFP buf_splitterG12ton164n259_splitterG12ton258n259_8_( clk_6 , buf_splitterG12ton164n259_splitterG12ton258n259_9 , 0 , buf_splitterG12ton164n259_splitterG12ton258n259_8 );
buf_AQFP buf_splitterG12ton164n259_splitterG12ton258n259_7_( clk_8 , buf_splitterG12ton164n259_splitterG12ton258n259_8 , 0 , buf_splitterG12ton164n259_splitterG12ton258n259_7 );
buf_AQFP buf_splitterG12ton164n259_splitterG12ton258n259_6_( clk_2 , buf_splitterG12ton164n259_splitterG12ton258n259_7 , 0 , buf_splitterG12ton164n259_splitterG12ton258n259_6 );
buf_AQFP buf_splitterG12ton164n259_splitterG12ton258n259_5_( clk_4 , buf_splitterG12ton164n259_splitterG12ton258n259_6 , 0 , buf_splitterG12ton164n259_splitterG12ton258n259_5 );
buf_AQFP buf_splitterG12ton164n259_splitterG12ton258n259_4_( clk_6 , buf_splitterG12ton164n259_splitterG12ton258n259_5 , 0 , buf_splitterG12ton164n259_splitterG12ton258n259_4 );
buf_AQFP buf_splitterG12ton164n259_splitterG12ton258n259_3_( clk_8 , buf_splitterG12ton164n259_splitterG12ton258n259_4 , 0 , buf_splitterG12ton164n259_splitterG12ton258n259_3 );
buf_AQFP buf_splitterG12ton164n259_splitterG12ton258n259_2_( clk_2 , buf_splitterG12ton164n259_splitterG12ton258n259_3 , 0 , buf_splitterG12ton164n259_splitterG12ton258n259_2 );
buf_AQFP buf_splitterG12ton164n259_splitterG12ton258n259_1_( clk_4 , buf_splitterG12ton164n259_splitterG12ton258n259_2 , 0 , buf_splitterG12ton164n259_splitterG12ton258n259_1 );
buf_AQFP buf_splitterG13ton79n262_splitterG13ton111n262_1_( clk_5 , splitterG13ton79n262 , 0 , buf_splitterG13ton79n262_splitterG13ton111n262_1 );
buf_AQFP buf_splitterG13ton111n262_splitterG13ton261n262_11_( clk_8 , splitterG13ton111n262 , 0 , buf_splitterG13ton111n262_splitterG13ton261n262_11 );
buf_AQFP buf_splitterG13ton111n262_splitterG13ton261n262_10_( clk_2 , buf_splitterG13ton111n262_splitterG13ton261n262_11 , 0 , buf_splitterG13ton111n262_splitterG13ton261n262_10 );
buf_AQFP buf_splitterG13ton111n262_splitterG13ton261n262_9_( clk_4 , buf_splitterG13ton111n262_splitterG13ton261n262_10 , 0 , buf_splitterG13ton111n262_splitterG13ton261n262_9 );
buf_AQFP buf_splitterG13ton111n262_splitterG13ton261n262_8_( clk_6 , buf_splitterG13ton111n262_splitterG13ton261n262_9 , 0 , buf_splitterG13ton111n262_splitterG13ton261n262_8 );
buf_AQFP buf_splitterG13ton111n262_splitterG13ton261n262_7_( clk_8 , buf_splitterG13ton111n262_splitterG13ton261n262_8 , 0 , buf_splitterG13ton111n262_splitterG13ton261n262_7 );
buf_AQFP buf_splitterG13ton111n262_splitterG13ton261n262_6_( clk_2 , buf_splitterG13ton111n262_splitterG13ton261n262_7 , 0 , buf_splitterG13ton111n262_splitterG13ton261n262_6 );
buf_AQFP buf_splitterG13ton111n262_splitterG13ton261n262_5_( clk_4 , buf_splitterG13ton111n262_splitterG13ton261n262_6 , 0 , buf_splitterG13ton111n262_splitterG13ton261n262_5 );
buf_AQFP buf_splitterG13ton111n262_splitterG13ton261n262_4_( clk_6 , buf_splitterG13ton111n262_splitterG13ton261n262_5 , 0 , buf_splitterG13ton111n262_splitterG13ton261n262_4 );
buf_AQFP buf_splitterG13ton111n262_splitterG13ton261n262_3_( clk_8 , buf_splitterG13ton111n262_splitterG13ton261n262_4 , 0 , buf_splitterG13ton111n262_splitterG13ton261n262_3 );
buf_AQFP buf_splitterG13ton111n262_splitterG13ton261n262_2_( clk_2 , buf_splitterG13ton111n262_splitterG13ton261n262_3 , 0 , buf_splitterG13ton111n262_splitterG13ton261n262_2 );
buf_AQFP buf_splitterG13ton111n262_splitterG13ton261n262_1_( clk_4 , buf_splitterG13ton111n262_splitterG13ton261n262_2 , 0 , buf_splitterG13ton111n262_splitterG13ton261n262_1 );
buf_AQFP buf_splitterG14ton103n265_splitterG14ton264n265_12_( clk_6 , splitterG14ton103n265 , 0 , buf_splitterG14ton103n265_splitterG14ton264n265_12 );
buf_AQFP buf_splitterG14ton103n265_splitterG14ton264n265_11_( clk_8 , buf_splitterG14ton103n265_splitterG14ton264n265_12 , 0 , buf_splitterG14ton103n265_splitterG14ton264n265_11 );
buf_AQFP buf_splitterG14ton103n265_splitterG14ton264n265_10_( clk_2 , buf_splitterG14ton103n265_splitterG14ton264n265_11 , 0 , buf_splitterG14ton103n265_splitterG14ton264n265_10 );
buf_AQFP buf_splitterG14ton103n265_splitterG14ton264n265_9_( clk_4 , buf_splitterG14ton103n265_splitterG14ton264n265_10 , 0 , buf_splitterG14ton103n265_splitterG14ton264n265_9 );
buf_AQFP buf_splitterG14ton103n265_splitterG14ton264n265_8_( clk_6 , buf_splitterG14ton103n265_splitterG14ton264n265_9 , 0 , buf_splitterG14ton103n265_splitterG14ton264n265_8 );
buf_AQFP buf_splitterG14ton103n265_splitterG14ton264n265_7_( clk_8 , buf_splitterG14ton103n265_splitterG14ton264n265_8 , 0 , buf_splitterG14ton103n265_splitterG14ton264n265_7 );
buf_AQFP buf_splitterG14ton103n265_splitterG14ton264n265_6_( clk_2 , buf_splitterG14ton103n265_splitterG14ton264n265_7 , 0 , buf_splitterG14ton103n265_splitterG14ton264n265_6 );
buf_AQFP buf_splitterG14ton103n265_splitterG14ton264n265_5_( clk_4 , buf_splitterG14ton103n265_splitterG14ton264n265_6 , 0 , buf_splitterG14ton103n265_splitterG14ton264n265_5 );
buf_AQFP buf_splitterG14ton103n265_splitterG14ton264n265_4_( clk_6 , buf_splitterG14ton103n265_splitterG14ton264n265_5 , 0 , buf_splitterG14ton103n265_splitterG14ton264n265_4 );
buf_AQFP buf_splitterG14ton103n265_splitterG14ton264n265_3_( clk_8 , buf_splitterG14ton103n265_splitterG14ton264n265_4 , 0 , buf_splitterG14ton103n265_splitterG14ton264n265_3 );
buf_AQFP buf_splitterG14ton103n265_splitterG14ton264n265_2_( clk_2 , buf_splitterG14ton103n265_splitterG14ton264n265_3 , 0 , buf_splitterG14ton103n265_splitterG14ton264n265_2 );
buf_AQFP buf_splitterG14ton103n265_splitterG14ton264n265_1_( clk_4 , buf_splitterG14ton103n265_splitterG14ton264n265_2 , 0 , buf_splitterG14ton103n265_splitterG14ton264n265_1 );
buf_AQFP buf_splitterG15ton135n227_splitterG15ton226n227_13_( clk_5 , splitterG15ton135n227 , 0 , buf_splitterG15ton135n227_splitterG15ton226n227_13 );
buf_AQFP buf_splitterG15ton135n227_splitterG15ton226n227_12_( clk_7 , buf_splitterG15ton135n227_splitterG15ton226n227_13 , 0 , buf_splitterG15ton135n227_splitterG15ton226n227_12 );
buf_AQFP buf_splitterG15ton135n227_splitterG15ton226n227_11_( clk_1 , buf_splitterG15ton135n227_splitterG15ton226n227_12 , 0 , buf_splitterG15ton135n227_splitterG15ton226n227_11 );
buf_AQFP buf_splitterG15ton135n227_splitterG15ton226n227_10_( clk_3 , buf_splitterG15ton135n227_splitterG15ton226n227_11 , 0 , buf_splitterG15ton135n227_splitterG15ton226n227_10 );
buf_AQFP buf_splitterG15ton135n227_splitterG15ton226n227_9_( clk_5 , buf_splitterG15ton135n227_splitterG15ton226n227_10 , 0 , buf_splitterG15ton135n227_splitterG15ton226n227_9 );
buf_AQFP buf_splitterG15ton135n227_splitterG15ton226n227_8_( clk_7 , buf_splitterG15ton135n227_splitterG15ton226n227_9 , 0 , buf_splitterG15ton135n227_splitterG15ton226n227_8 );
buf_AQFP buf_splitterG15ton135n227_splitterG15ton226n227_7_( clk_1 , buf_splitterG15ton135n227_splitterG15ton226n227_8 , 0 , buf_splitterG15ton135n227_splitterG15ton226n227_7 );
buf_AQFP buf_splitterG15ton135n227_splitterG15ton226n227_6_( clk_3 , buf_splitterG15ton135n227_splitterG15ton226n227_7 , 0 , buf_splitterG15ton135n227_splitterG15ton226n227_6 );
buf_AQFP buf_splitterG15ton135n227_splitterG15ton226n227_5_( clk_5 , buf_splitterG15ton135n227_splitterG15ton226n227_6 , 0 , buf_splitterG15ton135n227_splitterG15ton226n227_5 );
buf_AQFP buf_splitterG15ton135n227_splitterG15ton226n227_4_( clk_7 , buf_splitterG15ton135n227_splitterG15ton226n227_5 , 0 , buf_splitterG15ton135n227_splitterG15ton226n227_4 );
buf_AQFP buf_splitterG15ton135n227_splitterG15ton226n227_3_( clk_1 , buf_splitterG15ton135n227_splitterG15ton226n227_4 , 0 , buf_splitterG15ton135n227_splitterG15ton226n227_3 );
buf_AQFP buf_splitterG15ton135n227_splitterG15ton226n227_2_( clk_3 , buf_splitterG15ton135n227_splitterG15ton226n227_3 , 0 , buf_splitterG15ton135n227_splitterG15ton226n227_2 );
buf_AQFP buf_splitterG15ton135n227_splitterG15ton226n227_1_( clk_5 , buf_splitterG15ton135n227_splitterG15ton226n227_2 , 0 , buf_splitterG15ton135n227_splitterG15ton226n227_1 );
buf_AQFP buf_splitterG16ton64n230_n64_1_( clk_6 , splitterG16ton64n230 , 0 , buf_splitterG16ton64n230_n64_1 );
buf_AQFP buf_splitterG16ton65n230_splitterG16ton229n230_11_( clk_8 , splitterG16ton65n230 , 0 , buf_splitterG16ton65n230_splitterG16ton229n230_11 );
buf_AQFP buf_splitterG16ton65n230_splitterG16ton229n230_10_( clk_2 , buf_splitterG16ton65n230_splitterG16ton229n230_11 , 0 , buf_splitterG16ton65n230_splitterG16ton229n230_10 );
buf_AQFP buf_splitterG16ton65n230_splitterG16ton229n230_9_( clk_4 , buf_splitterG16ton65n230_splitterG16ton229n230_10 , 0 , buf_splitterG16ton65n230_splitterG16ton229n230_9 );
buf_AQFP buf_splitterG16ton65n230_splitterG16ton229n230_8_( clk_6 , buf_splitterG16ton65n230_splitterG16ton229n230_9 , 0 , buf_splitterG16ton65n230_splitterG16ton229n230_8 );
buf_AQFP buf_splitterG16ton65n230_splitterG16ton229n230_7_( clk_8 , buf_splitterG16ton65n230_splitterG16ton229n230_8 , 0 , buf_splitterG16ton65n230_splitterG16ton229n230_7 );
buf_AQFP buf_splitterG16ton65n230_splitterG16ton229n230_6_( clk_2 , buf_splitterG16ton65n230_splitterG16ton229n230_7 , 0 , buf_splitterG16ton65n230_splitterG16ton229n230_6 );
buf_AQFP buf_splitterG16ton65n230_splitterG16ton229n230_5_( clk_4 , buf_splitterG16ton65n230_splitterG16ton229n230_6 , 0 , buf_splitterG16ton65n230_splitterG16ton229n230_5 );
buf_AQFP buf_splitterG16ton65n230_splitterG16ton229n230_4_( clk_6 , buf_splitterG16ton65n230_splitterG16ton229n230_5 , 0 , buf_splitterG16ton65n230_splitterG16ton229n230_4 );
buf_AQFP buf_splitterG16ton65n230_splitterG16ton229n230_3_( clk_8 , buf_splitterG16ton65n230_splitterG16ton229n230_4 , 0 , buf_splitterG16ton65n230_splitterG16ton229n230_3 );
buf_AQFP buf_splitterG16ton65n230_splitterG16ton229n230_2_( clk_2 , buf_splitterG16ton65n230_splitterG16ton229n230_3 , 0 , buf_splitterG16ton65n230_splitterG16ton229n230_2 );
buf_AQFP buf_splitterG16ton65n230_splitterG16ton229n230_1_( clk_4 , buf_splitterG16ton65n230_splitterG16ton229n230_2 , 0 , buf_splitterG16ton65n230_splitterG16ton229n230_1 );
buf_AQFP buf_splitterfromG17_n74_1_( clk_6 , splitterfromG17 , 0 , buf_splitterfromG17_n74_1 );
buf_AQFP buf_splitterfromG18_n35_1_( clk_7 , splitterfromG18 , 0 , buf_splitterfromG18_n35_1 );
buf_AQFP buf_splitterfromG19_n128_1_( clk_6 , splitterfromG19 , 0 , buf_splitterfromG19_n128_1 );
buf_AQFP buf_splitterG2ton45n211_splitterG2ton146n211_2_( clk_5 , splitterG2ton45n211 , 0 , buf_splitterG2ton45n211_splitterG2ton146n211_2 );
buf_AQFP buf_splitterG2ton45n211_splitterG2ton146n211_1_( clk_7 , buf_splitterG2ton45n211_splitterG2ton146n211_2 , 0 , buf_splitterG2ton45n211_splitterG2ton146n211_1 );
buf_AQFP buf_splitterG2ton146n211_splitterG2ton210n211_10_( clk_2 , splitterG2ton146n211 , 0 , buf_splitterG2ton146n211_splitterG2ton210n211_10 );
buf_AQFP buf_splitterG2ton146n211_splitterG2ton210n211_9_( clk_4 , buf_splitterG2ton146n211_splitterG2ton210n211_10 , 0 , buf_splitterG2ton146n211_splitterG2ton210n211_9 );
buf_AQFP buf_splitterG2ton146n211_splitterG2ton210n211_8_( clk_6 , buf_splitterG2ton146n211_splitterG2ton210n211_9 , 0 , buf_splitterG2ton146n211_splitterG2ton210n211_8 );
buf_AQFP buf_splitterG2ton146n211_splitterG2ton210n211_7_( clk_8 , buf_splitterG2ton146n211_splitterG2ton210n211_8 , 0 , buf_splitterG2ton146n211_splitterG2ton210n211_7 );
buf_AQFP buf_splitterG2ton146n211_splitterG2ton210n211_6_( clk_2 , buf_splitterG2ton146n211_splitterG2ton210n211_7 , 0 , buf_splitterG2ton146n211_splitterG2ton210n211_6 );
buf_AQFP buf_splitterG2ton146n211_splitterG2ton210n211_5_( clk_4 , buf_splitterG2ton146n211_splitterG2ton210n211_6 , 0 , buf_splitterG2ton146n211_splitterG2ton210n211_5 );
buf_AQFP buf_splitterG2ton146n211_splitterG2ton210n211_4_( clk_6 , buf_splitterG2ton146n211_splitterG2ton210n211_5 , 0 , buf_splitterG2ton146n211_splitterG2ton210n211_4 );
buf_AQFP buf_splitterG2ton146n211_splitterG2ton210n211_3_( clk_8 , buf_splitterG2ton146n211_splitterG2ton210n211_4 , 0 , buf_splitterG2ton146n211_splitterG2ton210n211_3 );
buf_AQFP buf_splitterG2ton146n211_splitterG2ton210n211_2_( clk_2 , buf_splitterG2ton146n211_splitterG2ton210n211_3 , 0 , buf_splitterG2ton146n211_splitterG2ton210n211_2 );
buf_AQFP buf_splitterG2ton146n211_splitterG2ton210n211_1_( clk_4 , buf_splitterG2ton146n211_splitterG2ton210n211_2 , 0 , buf_splitterG2ton146n211_splitterG2ton210n211_1 );
buf_AQFP buf_splitterfromG20_n178_1_( clk_7 , splitterfromG20 , 0 , buf_splitterfromG20_n178_1 );
buf_AQFP buf_splitterG25ton193n281_n281_6_( clk_4 , splitterG25ton193n281 , 0 , buf_splitterG25ton193n281_n281_6 );
buf_AQFP buf_splitterG25ton193n281_n281_5_( clk_6 , buf_splitterG25ton193n281_n281_6 , 0 , buf_splitterG25ton193n281_n281_5 );
buf_AQFP buf_splitterG25ton193n281_n281_4_( clk_8 , buf_splitterG25ton193n281_n281_5 , 0 , buf_splitterG25ton193n281_n281_4 );
buf_AQFP buf_splitterG25ton193n281_n281_3_( clk_2 , buf_splitterG25ton193n281_n281_4 , 0 , buf_splitterG25ton193n281_n281_3 );
buf_AQFP buf_splitterG25ton193n281_n281_2_( clk_4 , buf_splitterG25ton193n281_n281_3 , 0 , buf_splitterG25ton193n281_n281_2 );
buf_AQFP buf_splitterG25ton193n281_n281_1_( clk_6 , buf_splitterG25ton193n281_n281_2 , 0 , buf_splitterG25ton193n281_n281_1 );
buf_AQFP buf_splitterG26ton100n320_n320_7_( clk_3 , splitterG26ton100n320 , 0 , buf_splitterG26ton100n320_n320_7 );
buf_AQFP buf_splitterG26ton100n320_n320_6_( clk_5 , buf_splitterG26ton100n320_n320_7 , 0 , buf_splitterG26ton100n320_n320_6 );
buf_AQFP buf_splitterG26ton100n320_n320_5_( clk_7 , buf_splitterG26ton100n320_n320_6 , 0 , buf_splitterG26ton100n320_n320_5 );
buf_AQFP buf_splitterG26ton100n320_n320_4_( clk_1 , buf_splitterG26ton100n320_n320_5 , 0 , buf_splitterG26ton100n320_n320_4 );
buf_AQFP buf_splitterG26ton100n320_n320_3_( clk_3 , buf_splitterG26ton100n320_n320_4 , 0 , buf_splitterG26ton100n320_n320_3 );
buf_AQFP buf_splitterG26ton100n320_n320_2_( clk_5 , buf_splitterG26ton100n320_n320_3 , 0 , buf_splitterG26ton100n320_n320_2 );
buf_AQFP buf_splitterG26ton100n320_n320_1_( clk_7 , buf_splitterG26ton100n320_n320_2 , 0 , buf_splitterG26ton100n320_n320_1 );
buf_AQFP buf_splitterG27ton153n287_n287_1_( clk_3 , splitterG27ton153n287 , 0 , buf_splitterG27ton153n287_n287_1 );
buf_AQFP buf_splitterG28ton173n291_n291_2_( clk_3 , splitterG28ton173n291 , 0 , buf_splitterG28ton173n291_n291_2 );
buf_AQFP buf_splitterG28ton173n291_n291_1_( clk_5 , buf_splitterG28ton173n291_n291_2 , 0 , buf_splitterG28ton173n291_n291_1 );
buf_AQFP buf_splitterfromG29_n199_1_( clk_6 , splitterfromG29 , 0 , buf_splitterfromG29_n199_1 );
buf_AQFP buf_splitterG3ton156n214_splitterG3ton213n214_12_( clk_7 , splitterG3ton156n214 , 0 , buf_splitterG3ton156n214_splitterG3ton213n214_12 );
buf_AQFP buf_splitterG3ton156n214_splitterG3ton213n214_11_( clk_1 , buf_splitterG3ton156n214_splitterG3ton213n214_12 , 0 , buf_splitterG3ton156n214_splitterG3ton213n214_11 );
buf_AQFP buf_splitterG3ton156n214_splitterG3ton213n214_10_( clk_3 , buf_splitterG3ton156n214_splitterG3ton213n214_11 , 0 , buf_splitterG3ton156n214_splitterG3ton213n214_10 );
buf_AQFP buf_splitterG3ton156n214_splitterG3ton213n214_9_( clk_5 , buf_splitterG3ton156n214_splitterG3ton213n214_10 , 0 , buf_splitterG3ton156n214_splitterG3ton213n214_9 );
buf_AQFP buf_splitterG3ton156n214_splitterG3ton213n214_8_( clk_7 , buf_splitterG3ton156n214_splitterG3ton213n214_9 , 0 , buf_splitterG3ton156n214_splitterG3ton213n214_8 );
buf_AQFP buf_splitterG3ton156n214_splitterG3ton213n214_7_( clk_1 , buf_splitterG3ton156n214_splitterG3ton213n214_8 , 0 , buf_splitterG3ton156n214_splitterG3ton213n214_7 );
buf_AQFP buf_splitterG3ton156n214_splitterG3ton213n214_6_( clk_3 , buf_splitterG3ton156n214_splitterG3ton213n214_7 , 0 , buf_splitterG3ton156n214_splitterG3ton213n214_6 );
buf_AQFP buf_splitterG3ton156n214_splitterG3ton213n214_5_( clk_5 , buf_splitterG3ton156n214_splitterG3ton213n214_6 , 0 , buf_splitterG3ton156n214_splitterG3ton213n214_5 );
buf_AQFP buf_splitterG3ton156n214_splitterG3ton213n214_4_( clk_7 , buf_splitterG3ton156n214_splitterG3ton213n214_5 , 0 , buf_splitterG3ton156n214_splitterG3ton213n214_4 );
buf_AQFP buf_splitterG3ton156n214_splitterG3ton213n214_3_( clk_1 , buf_splitterG3ton156n214_splitterG3ton213n214_4 , 0 , buf_splitterG3ton156n214_splitterG3ton213n214_3 );
buf_AQFP buf_splitterG3ton156n214_splitterG3ton213n214_2_( clk_3 , buf_splitterG3ton156n214_splitterG3ton213n214_3 , 0 , buf_splitterG3ton156n214_splitterG3ton213n214_2 );
buf_AQFP buf_splitterG3ton156n214_splitterG3ton213n214_1_( clk_5 , buf_splitterG3ton156n214_splitterG3ton213n214_2 , 0 , buf_splitterG3ton156n214_splitterG3ton213n214_1 );
buf_AQFP buf_splitterfromG30_n219_1_( clk_6 , splitterfromG30 , 0 , buf_splitterfromG30_n219_1 );
buf_AQFP buf_splitterG31ton127n282_splitterG31ton126n282_5_( clk_6 , splitterG31ton127n282 , 0 , buf_splitterG31ton127n282_splitterG31ton126n282_5 );
buf_AQFP buf_splitterG31ton127n282_splitterG31ton126n282_4_( clk_8 , buf_splitterG31ton127n282_splitterG31ton126n282_5 , 0 , buf_splitterG31ton127n282_splitterG31ton126n282_4 );
buf_AQFP buf_splitterG31ton127n282_splitterG31ton126n282_3_( clk_2 , buf_splitterG31ton127n282_splitterG31ton126n282_4 , 0 , buf_splitterG31ton127n282_splitterG31ton126n282_3 );
buf_AQFP buf_splitterG31ton127n282_splitterG31ton126n282_2_( clk_4 , buf_splitterG31ton127n282_splitterG31ton126n282_3 , 0 , buf_splitterG31ton127n282_splitterG31ton126n282_2 );
buf_AQFP buf_splitterG31ton127n282_splitterG31ton126n282_1_( clk_6 , buf_splitterG31ton127n282_splitterG31ton126n282_2 , 0 , buf_splitterG31ton127n282_splitterG31ton126n282_1 );
buf_AQFP buf_splitterG31ton291n282_splitterG31ton276n282_4_( clk_8 , splitterG31ton291n282 , 0 , buf_splitterG31ton291n282_splitterG31ton276n282_4 );
buf_AQFP buf_splitterG31ton291n282_splitterG31ton276n282_3_( clk_2 , buf_splitterG31ton291n282_splitterG31ton276n282_4 , 0 , buf_splitterG31ton291n282_splitterG31ton276n282_3 );
buf_AQFP buf_splitterG31ton291n282_splitterG31ton276n282_2_( clk_4 , buf_splitterG31ton291n282_splitterG31ton276n282_3 , 0 , buf_splitterG31ton291n282_splitterG31ton276n282_2 );
buf_AQFP buf_splitterG31ton291n282_splitterG31ton276n282_1_( clk_6 , buf_splitterG31ton291n282_splitterG31ton276n282_2 , 0 , buf_splitterG31ton291n282_splitterG31ton276n282_1 );
buf_AQFP buf_splitterfromG32_n268_9_( clk_8 , splitterfromG32 , 0 , buf_splitterfromG32_n268_9 );
buf_AQFP buf_splitterfromG32_n268_8_( clk_2 , buf_splitterfromG32_n268_9 , 0 , buf_splitterfromG32_n268_8 );
buf_AQFP buf_splitterfromG32_n268_7_( clk_4 , buf_splitterfromG32_n268_8 , 0 , buf_splitterfromG32_n268_7 );
buf_AQFP buf_splitterfromG32_n268_6_( clk_6 , buf_splitterfromG32_n268_7 , 0 , buf_splitterfromG32_n268_6 );
buf_AQFP buf_splitterfromG32_n268_5_( clk_8 , buf_splitterfromG32_n268_6 , 0 , buf_splitterfromG32_n268_5 );
buf_AQFP buf_splitterfromG32_n268_4_( clk_2 , buf_splitterfromG32_n268_5 , 0 , buf_splitterfromG32_n268_4 );
buf_AQFP buf_splitterfromG32_n268_3_( clk_4 , buf_splitterfromG32_n268_4 , 0 , buf_splitterfromG32_n268_3 );
buf_AQFP buf_splitterfromG32_n268_2_( clk_6 , buf_splitterfromG32_n268_3 , 0 , buf_splitterfromG32_n268_2 );
buf_AQFP buf_splitterfromG32_n268_1_( clk_8 , buf_splitterfromG32_n268_2 , 0 , buf_splitterfromG32_n268_1 );
buf_AQFP buf_splitterG33ton199n316_splitterG33ton203n316_3_( clk_1 , splitterG33ton199n316 , 0 , buf_splitterG33ton199n316_splitterG33ton203n316_3 );
buf_AQFP buf_splitterG33ton199n316_splitterG33ton203n316_2_( clk_3 , buf_splitterG33ton199n316_splitterG33ton203n316_3 , 0 , buf_splitterG33ton199n316_splitterG33ton203n316_2 );
buf_AQFP buf_splitterG33ton199n316_splitterG33ton203n316_1_( clk_5 , buf_splitterG33ton199n316_splitterG33ton203n316_2 , 0 , buf_splitterG33ton199n316_splitterG33ton203n316_1 );
buf_AQFP buf_splitterG33ton203n316_splitterG33ton273n316_7_( clk_1 , splitterG33ton203n316 , 0 , buf_splitterG33ton203n316_splitterG33ton273n316_7 );
buf_AQFP buf_splitterG33ton203n316_splitterG33ton273n316_6_( clk_3 , buf_splitterG33ton203n316_splitterG33ton273n316_7 , 0 , buf_splitterG33ton203n316_splitterG33ton273n316_6 );
buf_AQFP buf_splitterG33ton203n316_splitterG33ton273n316_5_( clk_5 , buf_splitterG33ton203n316_splitterG33ton273n316_6 , 0 , buf_splitterG33ton203n316_splitterG33ton273n316_5 );
buf_AQFP buf_splitterG33ton203n316_splitterG33ton273n316_4_( clk_7 , buf_splitterG33ton203n316_splitterG33ton273n316_5 , 0 , buf_splitterG33ton203n316_splitterG33ton273n316_4 );
buf_AQFP buf_splitterG33ton203n316_splitterG33ton273n316_3_( clk_1 , buf_splitterG33ton203n316_splitterG33ton273n316_4 , 0 , buf_splitterG33ton203n316_splitterG33ton273n316_3 );
buf_AQFP buf_splitterG33ton203n316_splitterG33ton273n316_2_( clk_3 , buf_splitterG33ton203n316_splitterG33ton273n316_3 , 0 , buf_splitterG33ton203n316_splitterG33ton273n316_2 );
buf_AQFP buf_splitterG33ton203n316_splitterG33ton273n316_1_( clk_5 , buf_splitterG33ton203n316_splitterG33ton273n316_2 , 0 , buf_splitterG33ton203n316_splitterG33ton273n316_1 );
buf_AQFP buf_splitterG4ton118n217_splitterG4ton216n217_11_( clk_8 , splitterG4ton118n217 , 0 , buf_splitterG4ton118n217_splitterG4ton216n217_11 );
buf_AQFP buf_splitterG4ton118n217_splitterG4ton216n217_10_( clk_2 , buf_splitterG4ton118n217_splitterG4ton216n217_11 , 0 , buf_splitterG4ton118n217_splitterG4ton216n217_10 );
buf_AQFP buf_splitterG4ton118n217_splitterG4ton216n217_9_( clk_4 , buf_splitterG4ton118n217_splitterG4ton216n217_10 , 0 , buf_splitterG4ton118n217_splitterG4ton216n217_9 );
buf_AQFP buf_splitterG4ton118n217_splitterG4ton216n217_8_( clk_6 , buf_splitterG4ton118n217_splitterG4ton216n217_9 , 0 , buf_splitterG4ton118n217_splitterG4ton216n217_8 );
buf_AQFP buf_splitterG4ton118n217_splitterG4ton216n217_7_( clk_8 , buf_splitterG4ton118n217_splitterG4ton216n217_8 , 0 , buf_splitterG4ton118n217_splitterG4ton216n217_7 );
buf_AQFP buf_splitterG4ton118n217_splitterG4ton216n217_6_( clk_2 , buf_splitterG4ton118n217_splitterG4ton216n217_7 , 0 , buf_splitterG4ton118n217_splitterG4ton216n217_6 );
buf_AQFP buf_splitterG4ton118n217_splitterG4ton216n217_5_( clk_4 , buf_splitterG4ton118n217_splitterG4ton216n217_6 , 0 , buf_splitterG4ton118n217_splitterG4ton216n217_5 );
buf_AQFP buf_splitterG4ton118n217_splitterG4ton216n217_4_( clk_6 , buf_splitterG4ton118n217_splitterG4ton216n217_5 , 0 , buf_splitterG4ton118n217_splitterG4ton216n217_4 );
buf_AQFP buf_splitterG4ton118n217_splitterG4ton216n217_3_( clk_8 , buf_splitterG4ton118n217_splitterG4ton216n217_4 , 0 , buf_splitterG4ton118n217_splitterG4ton216n217_3 );
buf_AQFP buf_splitterG4ton118n217_splitterG4ton216n217_2_( clk_2 , buf_splitterG4ton118n217_splitterG4ton216n217_3 , 0 , buf_splitterG4ton118n217_splitterG4ton216n217_2 );
buf_AQFP buf_splitterG4ton118n217_splitterG4ton216n217_1_( clk_4 , buf_splitterG4ton118n217_splitterG4ton216n217_2 , 0 , buf_splitterG4ton118n217_splitterG4ton216n217_1 );
buf_AQFP buf_splitterG5ton39n237_splitterG5ton236n237_10_( clk_8 , splitterG5ton39n237 , 0 , buf_splitterG5ton39n237_splitterG5ton236n237_10 );
buf_AQFP buf_splitterG5ton39n237_splitterG5ton236n237_9_( clk_2 , buf_splitterG5ton39n237_splitterG5ton236n237_10 , 0 , buf_splitterG5ton39n237_splitterG5ton236n237_9 );
buf_AQFP buf_splitterG5ton39n237_splitterG5ton236n237_8_( clk_4 , buf_splitterG5ton39n237_splitterG5ton236n237_9 , 0 , buf_splitterG5ton39n237_splitterG5ton236n237_8 );
buf_AQFP buf_splitterG5ton39n237_splitterG5ton236n237_7_( clk_6 , buf_splitterG5ton39n237_splitterG5ton236n237_8 , 0 , buf_splitterG5ton39n237_splitterG5ton236n237_7 );
buf_AQFP buf_splitterG5ton39n237_splitterG5ton236n237_6_( clk_8 , buf_splitterG5ton39n237_splitterG5ton236n237_7 , 0 , buf_splitterG5ton39n237_splitterG5ton236n237_6 );
buf_AQFP buf_splitterG5ton39n237_splitterG5ton236n237_5_( clk_2 , buf_splitterG5ton39n237_splitterG5ton236n237_6 , 0 , buf_splitterG5ton39n237_splitterG5ton236n237_5 );
buf_AQFP buf_splitterG5ton39n237_splitterG5ton236n237_4_( clk_4 , buf_splitterG5ton39n237_splitterG5ton236n237_5 , 0 , buf_splitterG5ton39n237_splitterG5ton236n237_4 );
buf_AQFP buf_splitterG5ton39n237_splitterG5ton236n237_3_( clk_6 , buf_splitterG5ton39n237_splitterG5ton236n237_4 , 0 , buf_splitterG5ton39n237_splitterG5ton236n237_3 );
buf_AQFP buf_splitterG5ton39n237_splitterG5ton236n237_2_( clk_8 , buf_splitterG5ton39n237_splitterG5ton236n237_3 , 0 , buf_splitterG5ton39n237_splitterG5ton236n237_2 );
buf_AQFP buf_splitterG5ton39n237_splitterG5ton236n237_1_( clk_2 , buf_splitterG5ton39n237_splitterG5ton236n237_2 , 0 , buf_splitterG5ton39n237_splitterG5ton236n237_1 );
buf_AQFP buf_splitterG6ton156n240_splitterG6ton239n240_11_( clk_7 , splitterG6ton156n240 , 0 , buf_splitterG6ton156n240_splitterG6ton239n240_11 );
buf_AQFP buf_splitterG6ton156n240_splitterG6ton239n240_10_( clk_1 , buf_splitterG6ton156n240_splitterG6ton239n240_11 , 0 , buf_splitterG6ton156n240_splitterG6ton239n240_10 );
buf_AQFP buf_splitterG6ton156n240_splitterG6ton239n240_9_( clk_3 , buf_splitterG6ton156n240_splitterG6ton239n240_10 , 0 , buf_splitterG6ton156n240_splitterG6ton239n240_9 );
buf_AQFP buf_splitterG6ton156n240_splitterG6ton239n240_8_( clk_5 , buf_splitterG6ton156n240_splitterG6ton239n240_9 , 0 , buf_splitterG6ton156n240_splitterG6ton239n240_8 );
buf_AQFP buf_splitterG6ton156n240_splitterG6ton239n240_7_( clk_7 , buf_splitterG6ton156n240_splitterG6ton239n240_8 , 0 , buf_splitterG6ton156n240_splitterG6ton239n240_7 );
buf_AQFP buf_splitterG6ton156n240_splitterG6ton239n240_6_( clk_1 , buf_splitterG6ton156n240_splitterG6ton239n240_7 , 0 , buf_splitterG6ton156n240_splitterG6ton239n240_6 );
buf_AQFP buf_splitterG6ton156n240_splitterG6ton239n240_5_( clk_3 , buf_splitterG6ton156n240_splitterG6ton239n240_6 , 0 , buf_splitterG6ton156n240_splitterG6ton239n240_5 );
buf_AQFP buf_splitterG6ton156n240_splitterG6ton239n240_4_( clk_5 , buf_splitterG6ton156n240_splitterG6ton239n240_5 , 0 , buf_splitterG6ton156n240_splitterG6ton239n240_4 );
buf_AQFP buf_splitterG6ton156n240_splitterG6ton239n240_3_( clk_7 , buf_splitterG6ton156n240_splitterG6ton239n240_4 , 0 , buf_splitterG6ton156n240_splitterG6ton239n240_3 );
buf_AQFP buf_splitterG6ton156n240_splitterG6ton239n240_2_( clk_1 , buf_splitterG6ton156n240_splitterG6ton239n240_3 , 0 , buf_splitterG6ton156n240_splitterG6ton239n240_2 );
buf_AQFP buf_splitterG6ton156n240_splitterG6ton239n240_1_( clk_3 , buf_splitterG6ton156n240_splitterG6ton239n240_2 , 0 , buf_splitterG6ton156n240_splitterG6ton239n240_1 );
buf_AQFP buf_splitterG7ton117n243_splitterG7ton242n243_11_( clk_7 , splitterG7ton117n243 , 0 , buf_splitterG7ton117n243_splitterG7ton242n243_11 );
buf_AQFP buf_splitterG7ton117n243_splitterG7ton242n243_10_( clk_1 , buf_splitterG7ton117n243_splitterG7ton242n243_11 , 0 , buf_splitterG7ton117n243_splitterG7ton242n243_10 );
buf_AQFP buf_splitterG7ton117n243_splitterG7ton242n243_9_( clk_3 , buf_splitterG7ton117n243_splitterG7ton242n243_10 , 0 , buf_splitterG7ton117n243_splitterG7ton242n243_9 );
buf_AQFP buf_splitterG7ton117n243_splitterG7ton242n243_8_( clk_5 , buf_splitterG7ton117n243_splitterG7ton242n243_9 , 0 , buf_splitterG7ton117n243_splitterG7ton242n243_8 );
buf_AQFP buf_splitterG7ton117n243_splitterG7ton242n243_7_( clk_7 , buf_splitterG7ton117n243_splitterG7ton242n243_8 , 0 , buf_splitterG7ton117n243_splitterG7ton242n243_7 );
buf_AQFP buf_splitterG7ton117n243_splitterG7ton242n243_6_( clk_1 , buf_splitterG7ton117n243_splitterG7ton242n243_7 , 0 , buf_splitterG7ton117n243_splitterG7ton242n243_6 );
buf_AQFP buf_splitterG7ton117n243_splitterG7ton242n243_5_( clk_3 , buf_splitterG7ton117n243_splitterG7ton242n243_6 , 0 , buf_splitterG7ton117n243_splitterG7ton242n243_5 );
buf_AQFP buf_splitterG7ton117n243_splitterG7ton242n243_4_( clk_5 , buf_splitterG7ton117n243_splitterG7ton242n243_5 , 0 , buf_splitterG7ton117n243_splitterG7ton242n243_4 );
buf_AQFP buf_splitterG7ton117n243_splitterG7ton242n243_3_( clk_7 , buf_splitterG7ton117n243_splitterG7ton242n243_4 , 0 , buf_splitterG7ton117n243_splitterG7ton242n243_3 );
buf_AQFP buf_splitterG7ton117n243_splitterG7ton242n243_2_( clk_1 , buf_splitterG7ton117n243_splitterG7ton242n243_3 , 0 , buf_splitterG7ton117n243_splitterG7ton242n243_2 );
buf_AQFP buf_splitterG7ton117n243_splitterG7ton242n243_1_( clk_3 , buf_splitterG7ton117n243_splitterG7ton242n243_2 , 0 , buf_splitterG7ton117n243_splitterG7ton242n243_1 );
buf_AQFP buf_splitterG8ton159n246_splitterG8ton245n246_10_( clk_1 , splitterG8ton159n246 , 0 , buf_splitterG8ton159n246_splitterG8ton245n246_10 );
buf_AQFP buf_splitterG8ton159n246_splitterG8ton245n246_9_( clk_3 , buf_splitterG8ton159n246_splitterG8ton245n246_10 , 0 , buf_splitterG8ton159n246_splitterG8ton245n246_9 );
buf_AQFP buf_splitterG8ton159n246_splitterG8ton245n246_8_( clk_5 , buf_splitterG8ton159n246_splitterG8ton245n246_9 , 0 , buf_splitterG8ton159n246_splitterG8ton245n246_8 );
buf_AQFP buf_splitterG8ton159n246_splitterG8ton245n246_7_( clk_7 , buf_splitterG8ton159n246_splitterG8ton245n246_8 , 0 , buf_splitterG8ton159n246_splitterG8ton245n246_7 );
buf_AQFP buf_splitterG8ton159n246_splitterG8ton245n246_6_( clk_1 , buf_splitterG8ton159n246_splitterG8ton245n246_7 , 0 , buf_splitterG8ton159n246_splitterG8ton245n246_6 );
buf_AQFP buf_splitterG8ton159n246_splitterG8ton245n246_5_( clk_3 , buf_splitterG8ton159n246_splitterG8ton245n246_6 , 0 , buf_splitterG8ton159n246_splitterG8ton245n246_5 );
buf_AQFP buf_splitterG8ton159n246_splitterG8ton245n246_4_( clk_5 , buf_splitterG8ton159n246_splitterG8ton245n246_5 , 0 , buf_splitterG8ton159n246_splitterG8ton245n246_4 );
buf_AQFP buf_splitterG8ton159n246_splitterG8ton245n246_3_( clk_7 , buf_splitterG8ton159n246_splitterG8ton245n246_4 , 0 , buf_splitterG8ton159n246_splitterG8ton245n246_3 );
buf_AQFP buf_splitterG8ton159n246_splitterG8ton245n246_2_( clk_1 , buf_splitterG8ton159n246_splitterG8ton245n246_3 , 0 , buf_splitterG8ton159n246_splitterG8ton245n246_2 );
buf_AQFP buf_splitterG8ton159n246_splitterG8ton245n246_1_( clk_3 , buf_splitterG8ton159n246_splitterG8ton245n246_2 , 0 , buf_splitterG8ton159n246_splitterG8ton245n246_1 );
buf_AQFP buf_splitterG9ton103n250_splitterG9ton58n250_1_( clk_5 , splitterG9ton103n250 , 0 , buf_splitterG9ton103n250_splitterG9ton58n250_1 );
buf_AQFP buf_splitterG9ton58n250_splitterG9ton249n250_10_( clk_1 , splitterG9ton58n250 , 0 , buf_splitterG9ton58n250_splitterG9ton249n250_10 );
buf_AQFP buf_splitterG9ton58n250_splitterG9ton249n250_9_( clk_3 , buf_splitterG9ton58n250_splitterG9ton249n250_10 , 0 , buf_splitterG9ton58n250_splitterG9ton249n250_9 );
buf_AQFP buf_splitterG9ton58n250_splitterG9ton249n250_8_( clk_5 , buf_splitterG9ton58n250_splitterG9ton249n250_9 , 0 , buf_splitterG9ton58n250_splitterG9ton249n250_8 );
buf_AQFP buf_splitterG9ton58n250_splitterG9ton249n250_7_( clk_7 , buf_splitterG9ton58n250_splitterG9ton249n250_8 , 0 , buf_splitterG9ton58n250_splitterG9ton249n250_7 );
buf_AQFP buf_splitterG9ton58n250_splitterG9ton249n250_6_( clk_1 , buf_splitterG9ton58n250_splitterG9ton249n250_7 , 0 , buf_splitterG9ton58n250_splitterG9ton249n250_6 );
buf_AQFP buf_splitterG9ton58n250_splitterG9ton249n250_5_( clk_3 , buf_splitterG9ton58n250_splitterG9ton249n250_6 , 0 , buf_splitterG9ton58n250_splitterG9ton249n250_5 );
buf_AQFP buf_splitterG9ton58n250_splitterG9ton249n250_4_( clk_5 , buf_splitterG9ton58n250_splitterG9ton249n250_5 , 0 , buf_splitterG9ton58n250_splitterG9ton249n250_4 );
buf_AQFP buf_splitterG9ton58n250_splitterG9ton249n250_3_( clk_7 , buf_splitterG9ton58n250_splitterG9ton249n250_4 , 0 , buf_splitterG9ton58n250_splitterG9ton249n250_3 );
buf_AQFP buf_splitterG9ton58n250_splitterG9ton249n250_2_( clk_1 , buf_splitterG9ton58n250_splitterG9ton249n250_3 , 0 , buf_splitterG9ton58n250_splitterG9ton249n250_2 );
buf_AQFP buf_splitterG9ton58n250_splitterG9ton249n250_1_( clk_3 , buf_splitterG9ton58n250_splitterG9ton249n250_2 , 0 , buf_splitterG9ton58n250_splitterG9ton249n250_1 );
buf_AQFP buf_splittern35ton78n252_n252_1_( clk_8 , splittern35ton78n252 , 0 , buf_splittern35ton78n252_n252_1 );
buf_AQFP buf_splitterfromn72_n277_8_( clk_4 , splitterfromn72 , 0 , buf_splitterfromn72_n277_8 );
buf_AQFP buf_splitterfromn72_n277_7_( clk_6 , buf_splitterfromn72_n277_8 , 0 , buf_splitterfromn72_n277_7 );
buf_AQFP buf_splitterfromn72_n277_6_( clk_8 , buf_splitterfromn72_n277_7 , 0 , buf_splitterfromn72_n277_6 );
buf_AQFP buf_splitterfromn72_n277_5_( clk_2 , buf_splitterfromn72_n277_6 , 0 , buf_splitterfromn72_n277_5 );
buf_AQFP buf_splitterfromn72_n277_4_( clk_4 , buf_splitterfromn72_n277_5 , 0 , buf_splitterfromn72_n277_4 );
buf_AQFP buf_splitterfromn72_n277_3_( clk_6 , buf_splitterfromn72_n277_4 , 0 , buf_splitterfromn72_n277_3 );
buf_AQFP buf_splitterfromn72_n277_2_( clk_8 , buf_splitterfromn72_n277_3 , 0 , buf_splitterfromn72_n277_2 );
buf_AQFP buf_splitterfromn72_n277_1_( clk_2 , buf_splitterfromn72_n277_2 , 0 , buf_splitterfromn72_n277_1 );
buf_AQFP buf_splittern73ton75n278_n278_6_( clk_6 , splittern73ton75n278 , 0 , buf_splittern73ton75n278_n278_6 );
buf_AQFP buf_splittern73ton75n278_n278_5_( clk_8 , buf_splittern73ton75n278_n278_6 , 0 , buf_splittern73ton75n278_n278_5 );
buf_AQFP buf_splittern73ton75n278_n278_4_( clk_2 , buf_splittern73ton75n278_n278_5 , 0 , buf_splittern73ton75n278_n278_4 );
buf_AQFP buf_splittern73ton75n278_n278_3_( clk_4 , buf_splittern73ton75n278_n278_4 , 0 , buf_splittern73ton75n278_n278_3 );
buf_AQFP buf_splittern73ton75n278_n278_2_( clk_6 , buf_splittern73ton75n278_n278_3 , 0 , buf_splittern73ton75n278_n278_2 );
buf_AQFP buf_splittern73ton75n278_n278_1_( clk_8 , buf_splittern73ton75n278_n278_2 , 0 , buf_splittern73ton75n278_n278_1 );
buf_AQFP buf_splittern74ton75n275_n275_6_( clk_5 , splittern74ton75n275 , 0 , buf_splittern74ton75n275_n275_6 );
buf_AQFP buf_splittern74ton75n275_n275_5_( clk_7 , buf_splittern74ton75n275_n275_6 , 0 , buf_splittern74ton75n275_n275_5 );
buf_AQFP buf_splittern74ton75n275_n275_4_( clk_1 , buf_splittern74ton75n275_n275_5 , 0 , buf_splittern74ton75n275_n275_4 );
buf_AQFP buf_splittern74ton75n275_n275_3_( clk_3 , buf_splittern74ton75n275_n275_4 , 0 , buf_splittern74ton75n275_n275_3 );
buf_AQFP buf_splittern74ton75n275_n275_2_( clk_5 , buf_splittern74ton75n275_n275_3 , 0 , buf_splittern74ton75n275_n275_2 );
buf_AQFP buf_splittern74ton75n275_n275_1_( clk_7 , buf_splittern74ton75n275_n275_2 , 0 , buf_splittern74ton75n275_n275_1 );
buf_AQFP buf_splittern77ton271n253_n253_1_( clk_1 , splittern77ton271n253 , 0 , buf_splittern77ton271n253_n253_1 );
buf_AQFP buf_splitterfromn98_n321_7_( clk_2 , splitterfromn98 , 0 , buf_splitterfromn98_n321_7 );
buf_AQFP buf_splitterfromn98_n321_6_( clk_4 , buf_splitterfromn98_n321_7 , 0 , buf_splitterfromn98_n321_6 );
buf_AQFP buf_splitterfromn98_n321_5_( clk_6 , buf_splitterfromn98_n321_6 , 0 , buf_splitterfromn98_n321_5 );
buf_AQFP buf_splitterfromn98_n321_4_( clk_8 , buf_splitterfromn98_n321_5 , 0 , buf_splitterfromn98_n321_4 );
buf_AQFP buf_splitterfromn98_n321_3_( clk_2 , buf_splitterfromn98_n321_4 , 0 , buf_splitterfromn98_n321_3 );
buf_AQFP buf_splitterfromn98_n321_2_( clk_4 , buf_splitterfromn98_n321_3 , 0 , buf_splitterfromn98_n321_2 );
buf_AQFP buf_splitterfromn98_n321_1_( clk_6 , buf_splitterfromn98_n321_2 , 0 , buf_splitterfromn98_n321_1 );
buf_AQFP buf_splittern105ton106n309_splittern105ton308n309_2_( clk_1 , splittern105ton106n309 , 0 , buf_splittern105ton106n309_splittern105ton308n309_2 );
buf_AQFP buf_splittern105ton106n309_splittern105ton308n309_1_( clk_3 , buf_splittern105ton106n309_splittern105ton308n309_2 , 0 , buf_splittern105ton106n309_splittern105ton308n309_1 );
buf_AQFP buf_splitterfromn125_n297_8_( clk_2 , splitterfromn125 , 0 , buf_splitterfromn125_n297_8 );
buf_AQFP buf_splitterfromn125_n297_7_( clk_4 , buf_splitterfromn125_n297_8 , 0 , buf_splitterfromn125_n297_7 );
buf_AQFP buf_splitterfromn125_n297_6_( clk_6 , buf_splitterfromn125_n297_7 , 0 , buf_splitterfromn125_n297_6 );
buf_AQFP buf_splitterfromn125_n297_5_( clk_8 , buf_splitterfromn125_n297_6 , 0 , buf_splitterfromn125_n297_5 );
buf_AQFP buf_splitterfromn125_n297_4_( clk_2 , buf_splitterfromn125_n297_5 , 0 , buf_splitterfromn125_n297_4 );
buf_AQFP buf_splitterfromn125_n297_3_( clk_4 , buf_splitterfromn125_n297_4 , 0 , buf_splitterfromn125_n297_3 );
buf_AQFP buf_splitterfromn125_n297_2_( clk_6 , buf_splitterfromn125_n297_3 , 0 , buf_splitterfromn125_n297_2 );
buf_AQFP buf_splitterfromn125_n297_1_( clk_8 , buf_splitterfromn125_n297_2 , 0 , buf_splitterfromn125_n297_1 );
buf_AQFP buf_splittern128ton129n295_n295_2_( clk_3 , splittern128ton129n295 , 0 , buf_splittern128ton129n295_n295_2 );
buf_AQFP buf_splittern128ton129n295_n295_1_( clk_5 , buf_splittern128ton129n295_n295_2 , 0 , buf_splittern128ton129n295_n295_1 );
buf_AQFP buf_splitterfromn151_n289_8_( clk_2 , splitterfromn151 , 0 , buf_splitterfromn151_n289_8 );
buf_AQFP buf_splitterfromn151_n289_7_( clk_4 , buf_splitterfromn151_n289_8 , 0 , buf_splitterfromn151_n289_7 );
buf_AQFP buf_splitterfromn151_n289_6_( clk_6 , buf_splitterfromn151_n289_7 , 0 , buf_splitterfromn151_n289_6 );
buf_AQFP buf_splitterfromn151_n289_5_( clk_8 , buf_splitterfromn151_n289_6 , 0 , buf_splitterfromn151_n289_5 );
buf_AQFP buf_splitterfromn151_n289_4_( clk_2 , buf_splitterfromn151_n289_5 , 0 , buf_splitterfromn151_n289_4 );
buf_AQFP buf_splitterfromn151_n289_3_( clk_4 , buf_splitterfromn151_n289_4 , 0 , buf_splitterfromn151_n289_3 );
buf_AQFP buf_splitterfromn151_n289_2_( clk_6 , buf_splitterfromn151_n289_3 , 0 , buf_splitterfromn151_n289_2 );
buf_AQFP buf_splitterfromn151_n289_1_( clk_8 , buf_splitterfromn151_n289_2 , 0 , buf_splitterfromn151_n289_1 );
buf_AQFP buf_splitterfromn171_n293_8_( clk_2 , splitterfromn171 , 0 , buf_splitterfromn171_n293_8 );
buf_AQFP buf_splitterfromn171_n293_7_( clk_4 , buf_splitterfromn171_n293_8 , 0 , buf_splitterfromn171_n293_7 );
buf_AQFP buf_splitterfromn171_n293_6_( clk_6 , buf_splitterfromn171_n293_7 , 0 , buf_splitterfromn171_n293_6 );
buf_AQFP buf_splitterfromn171_n293_5_( clk_8 , buf_splitterfromn171_n293_6 , 0 , buf_splitterfromn171_n293_5 );
buf_AQFP buf_splitterfromn171_n293_4_( clk_2 , buf_splitterfromn171_n293_5 , 0 , buf_splitterfromn171_n293_4 );
buf_AQFP buf_splitterfromn171_n293_3_( clk_4 , buf_splitterfromn171_n293_4 , 0 , buf_splitterfromn171_n293_3 );
buf_AQFP buf_splitterfromn171_n293_2_( clk_6 , buf_splitterfromn171_n293_3 , 0 , buf_splitterfromn171_n293_2 );
buf_AQFP buf_splitterfromn171_n293_1_( clk_8 , buf_splitterfromn171_n293_2 , 0 , buf_splitterfromn171_n293_1 );
buf_AQFP buf_splittern177ton197n272_n272_1_( clk_1 , splittern177ton197n272 , 0 , buf_splittern177ton197n272_n272_1 );
buf_AQFP buf_splitterfromn191_n283_8_( clk_3 , splitterfromn191 , 0 , buf_splitterfromn191_n283_8 );
buf_AQFP buf_splitterfromn191_n283_7_( clk_5 , buf_splitterfromn191_n283_8 , 0 , buf_splitterfromn191_n283_7 );
buf_AQFP buf_splitterfromn191_n283_6_( clk_7 , buf_splitterfromn191_n283_7 , 0 , buf_splitterfromn191_n283_6 );
buf_AQFP buf_splitterfromn191_n283_5_( clk_1 , buf_splitterfromn191_n283_6 , 0 , buf_splitterfromn191_n283_5 );
buf_AQFP buf_splitterfromn191_n283_4_( clk_3 , buf_splitterfromn191_n283_5 , 0 , buf_splitterfromn191_n283_4 );
buf_AQFP buf_splitterfromn191_n283_3_( clk_5 , buf_splitterfromn191_n283_4 , 0 , buf_splitterfromn191_n283_3 );
buf_AQFP buf_splitterfromn191_n283_2_( clk_7 , buf_splitterfromn191_n283_3 , 0 , buf_splitterfromn191_n283_2 );
buf_AQFP buf_splitterfromn191_n283_1_( clk_1 , buf_splitterfromn191_n283_2 , 0 , buf_splitterfromn191_n283_1 );
buf_AQFP buf_splittern192ton193n284_n284_7_( clk_5 , splittern192ton193n284 , 0 , buf_splittern192ton193n284_n284_7 );
buf_AQFP buf_splittern192ton193n284_n284_6_( clk_7 , buf_splittern192ton193n284_n284_7 , 0 , buf_splittern192ton193n284_n284_6 );
buf_AQFP buf_splittern192ton193n284_n284_5_( clk_1 , buf_splittern192ton193n284_n284_6 , 0 , buf_splittern192ton193n284_n284_5 );
buf_AQFP buf_splittern192ton193n284_n284_4_( clk_3 , buf_splittern192ton193n284_n284_5 , 0 , buf_splittern192ton193n284_n284_4 );
buf_AQFP buf_splittern192ton193n284_n284_3_( clk_5 , buf_splittern192ton193n284_n284_4 , 0 , buf_splittern192ton193n284_n284_3 );
buf_AQFP buf_splittern192ton193n284_n284_2_( clk_7 , buf_splittern192ton193n284_n284_3 , 0 , buf_splittern192ton193n284_n284_2 );
buf_AQFP buf_splittern192ton193n284_n284_1_( clk_1 , buf_splittern192ton193n284_n284_2 , 0 , buf_splittern192ton193n284_n284_1 );
buf_AQFP buf_splitterfromn199_n202_2_( clk_1 , splitterfromn199 , 0 , buf_splitterfromn199_n202_2 );
buf_AQFP buf_splitterfromn199_n202_1_( clk_3 , buf_splitterfromn199_n202_2 , 0 , buf_splitterfromn199_n202_1 );
buf_AQFP buf_splittern203ton204n298_splittern203ton321n298_5_( clk_4 , splittern203ton204n298 , 0 , buf_splittern203ton204n298_splittern203ton321n298_5 );
buf_AQFP buf_splittern203ton204n298_splittern203ton321n298_4_( clk_6 , buf_splittern203ton204n298_splittern203ton321n298_5 , 0 , buf_splittern203ton204n298_splittern203ton321n298_4 );
buf_AQFP buf_splittern203ton204n298_splittern203ton321n298_3_( clk_8 , buf_splittern203ton204n298_splittern203ton321n298_4 , 0 , buf_splittern203ton204n298_splittern203ton321n298_3 );
buf_AQFP buf_splittern203ton204n298_splittern203ton321n298_2_( clk_2 , buf_splittern203ton204n298_splittern203ton321n298_3 , 0 , buf_splittern203ton204n298_splittern203ton321n298_2 );
buf_AQFP buf_splittern203ton204n298_splittern203ton321n298_1_( clk_4 , buf_splittern203ton204n298_splittern203ton321n298_2 , 0 , buf_splittern203ton204n298_splittern203ton321n298_1 );
buf_AQFP buf_splittern203ton279n298_n279_1_( clk_1 , splittern203ton279n298 , 0 , buf_splittern203ton279n298_n279_1 );
buf_AQFP buf_splitterfromn219_n220_3_( clk_8 , splitterfromn219 , 0 , buf_splitterfromn219_n220_3 );
buf_AQFP buf_splitterfromn219_n220_2_( clk_2 , buf_splitterfromn219_n220_3 , 0 , buf_splitterfromn219_n220_2 );
buf_AQFP buf_splitterfromn219_n220_1_( clk_4 , buf_splitterfromn219_n220_2 , 0 , buf_splitterfromn219_n220_1 );
splitter_AQFP splitterG1ton48n208_( clk_4 , buf_G1_splitterG1ton48n208_1 , 0 , splitterG1ton48n208 );
splitter_AQFP splitterG1ton49n208_( clk_6 , splitterG1ton48n208 , 0 , splitterG1ton49n208 );
splitter_AQFP splitterG1ton207n208_( clk_6 , buf_splitterG1ton49n208_splitterG1ton207n208_1 , 0 , splitterG1ton207n208 );
splitter_AQFP splitterG10ton61n224_( clk_3 , G10 , 0 , splitterG10ton61n224 );
splitter_AQFP splitterG10ton120n224_( clk_8 , buf_splitterG10ton61n224_splitterG10ton120n224_1 , 0 , splitterG10ton120n224 );
splitter_AQFP splitterG10ton223n224_( clk_5 , buf_splitterG10ton120n224_splitterG10ton223n224_1 , 0 , splitterG10ton223n224 );
splitter_AQFP splitterG11ton134n256_( clk_2 , G11 , 0 , splitterG11ton134n256 );
splitter_AQFP splitterG11ton135n256_( clk_3 , splitterG11ton134n256 , 0 , splitterG11ton135n256 );
splitter_AQFP splitterG11ton255n256_( clk_5 , buf_splitterG11ton135n256_splitterG11ton255n256_1 , 0 , splitterG11ton255n256 );
splitter_AQFP splitterG12ton163n259_( clk_4 , buf_G12_splitterG12ton163n259_1 , 0 , splitterG12ton163n259 );
splitter_AQFP splitterG12ton164n259_( clk_6 , splitterG12ton163n259 , 0 , splitterG12ton164n259 );
splitter_AQFP splitterG12ton258n259_( clk_5 , buf_splitterG12ton164n259_splitterG12ton258n259_1 , 0 , splitterG12ton258n259 );
splitter_AQFP splitterG13ton79n262_( clk_3 , G13 , 0 , splitterG13ton79n262 );
splitter_AQFP splitterG13ton111n262_( clk_6 , buf_splitterG13ton79n262_splitterG13ton111n262_1 , 0 , splitterG13ton111n262 );
splitter_AQFP splitterG13ton261n262_( clk_5 , buf_splitterG13ton111n262_splitterG13ton261n262_1 , 0 , splitterG13ton261n262 );
splitter_AQFP splitterG14ton180n265_( clk_2 , G14 , 0 , splitterG14ton180n265 );
splitter_AQFP splitterG14ton103n265_( clk_4 , splitterG14ton180n265 , 0 , splitterG14ton103n265 );
splitter_AQFP splitterG14ton264n265_( clk_5 , buf_splitterG14ton103n265_splitterG14ton264n265_1 , 0 , splitterG14ton264n265 );
splitter_AQFP splitterG15ton134n227_( clk_2 , G15 , 0 , splitterG15ton134n227 );
splitter_AQFP splitterG15ton135n227_( clk_3 , splitterG15ton134n227 , 0 , splitterG15ton135n227 );
splitter_AQFP splitterG15ton226n227_( clk_6 , buf_splitterG15ton135n227_splitterG15ton226n227_1 , 0 , splitterG15ton226n227 );
splitter_AQFP splitterG16ton64n230_( clk_4 , buf_G16_splitterG16ton64n230_1 , 0 , splitterG16ton64n230 );
splitter_AQFP splitterG16ton65n230_( clk_6 , splitterG16ton64n230 , 0 , splitterG16ton65n230 );
splitter_AQFP splitterG16ton229n230_( clk_6 , buf_splitterG16ton65n230_splitterG16ton229n230_1 , 0 , splitterG16ton229n230 );
splitter_AQFP splitterfromG17_( clk_4 , buf_G17_splitterfromG17_1 , 0 , splitterfromG17 );
splitter_AQFP splitterfromG18_( clk_5 , buf_G18_splitterfromG18_1 , 0 , splitterfromG18 );
splitter_AQFP splitterfromG19_( clk_4 , buf_G19_splitterfromG19_1 , 0 , splitterfromG19 );
splitter_AQFP splitterG2ton45n211_( clk_3 , G2 , 0 , splitterG2ton45n211 );
splitter_AQFP splitterG2ton146n211_( clk_8 , buf_splitterG2ton45n211_splitterG2ton146n211_1 , 0 , splitterG2ton146n211 );
splitter_AQFP splitterG2ton210n211_( clk_6 , buf_splitterG2ton146n211_splitterG2ton210n211_1 , 0 , splitterG2ton210n211 );
splitter_AQFP splitterfromG20_( clk_5 , buf_G20_splitterfromG20_1 , 0 , splitterfromG20 );
splitter_AQFP splitterfromG21_( clk_4 , buf_G21_splitterfromG21_1 , 0 , splitterfromG21 );
splitter_AQFP splitterfromG22_( clk_4 , buf_G22_splitterfromG22_1 , 0 , splitterfromG22 );
splitter_AQFP splitterG23ton109n200_( clk_3 , G23 , 0 , splitterG23ton109n200 );
splitter_AQFP splitterG23ton127n200_( clk_5 , splitterG23ton109n200 , 0 , splitterG23ton127n200 );
splitter_AQFP splitterG24ton88n200_( clk_3 , G24 , 0 , splitterG24ton88n200 );
splitter_AQFP splitterG24ton34n200_( clk_5 , splitterG24ton88n200 , 0 , splitterG24ton34n200 );
splitter_AQFP splitterG25ton193n281_( clk_2 , buf_G25_splitterG25ton193n281_1 , 0 , splitterG25ton193n281 );
splitter_AQFP splitterG26ton100n320_( clk_1 , buf_G26_splitterG26ton100n320_1 , 0 , splitterG26ton100n320 );
splitter_AQFP splitterG27ton153n287_( clk_1 , buf_G27_splitterG27ton153n287_1 , 0 , splitterG27ton153n287 );
splitter_AQFP splitterG28ton173n291_( clk_1 , buf_G28_splitterG28ton173n291_1 , 0 , splitterG28ton173n291 );
splitter_AQFP splitterfromG29_( clk_4 , buf_G29_splitterfromG29_1 , 0 , splitterfromG29 );
splitter_AQFP splitterG3ton45n214_( clk_3 , G3 , 0 , splitterG3ton45n214 );
splitter_AQFP splitterG3ton156n214_( clk_5 , splitterG3ton45n214 , 0 , splitterG3ton156n214 );
splitter_AQFP splitterG3ton213n214_( clk_6 , buf_splitterG3ton156n214_splitterG3ton213n214_1 , 0 , splitterG3ton213n214 );
splitter_AQFP splitterfromG30_( clk_4 , buf_G30_splitterfromG30_1 , 0 , splitterfromG30 );
splitter_AQFP splitterG31ton127n282_( clk_4 , buf_G31_splitterG31ton127n282_1 , 0 , splitterG31ton127n282 );
splitter_AQFP splitterG31ton126n282_( clk_7 , buf_splitterG31ton127n282_splitterG31ton126n282_1 , 0 , splitterG31ton126n282 );
splitter_AQFP splitterG31ton172n282_( clk_8 , splitterG31ton126n282 , 0 , splitterG31ton172n282 );
splitter_AQFP splitterG31ton201n282_( clk_2 , splitterG31ton172n282 , 0 , splitterG31ton201n282 );
splitter_AQFP splitterG31ton287n282_( clk_4 , splitterG31ton201n282 , 0 , splitterG31ton287n282 );
splitter_AQFP splitterG31ton291n282_( clk_6 , splitterG31ton287n282 , 0 , splitterG31ton291n282 );
splitter_AQFP splitterG31ton276n282_( clk_8 , buf_splitterG31ton291n282_splitterG31ton276n282_1 , 0 , splitterG31ton276n282 );
splitter_AQFP splitterfromG32_( clk_6 , buf_G32_splitterfromG32_1 , 0 , splitterfromG32 );
splitter_AQFP splitterG33ton109n316_( clk_3 , G33 , 0 , splitterG33ton109n316 );
splitter_AQFP splitterG33ton179n316_( clk_5 , splitterG33ton109n316 , 0 , splitterG33ton179n316 );
splitter_AQFP splitterG33ton199n316_( clk_7 , splitterG33ton179n316 , 0 , splitterG33ton199n316 );
splitter_AQFP splitterG33ton203n316_( clk_7 , buf_splitterG33ton199n316_splitterG33ton203n316_1 , 0 , splitterG33ton203n316 );
splitter_AQFP splitterG33ton273n316_( clk_6 , buf_splitterG33ton203n316_splitterG33ton273n316_1 , 0 , splitterG33ton273n316 );
splitter_AQFP splitterG4ton180n217_( clk_2 , G4 , 0 , splitterG4ton180n217 );
splitter_AQFP splitterG4ton181n217_( clk_4 , splitterG4ton180n217 , 0 , splitterG4ton181n217 );
splitter_AQFP splitterG4ton118n217_( clk_6 , splitterG4ton181n217 , 0 , splitterG4ton118n217 );
splitter_AQFP splitterG4ton216n217_( clk_6 , buf_splitterG4ton118n217_splitterG4ton216n217_1 , 0 , splitterG4ton216n217 );
splitter_AQFP splitterG5ton143n237_( clk_4 , buf_G5_splitterG5ton143n237_1 , 0 , splitterG5ton143n237 );
splitter_AQFP splitterG5ton39n237_( clk_6 , splitterG5ton143n237 , 0 , splitterG5ton39n237 );
splitter_AQFP splitterG5ton236n237_( clk_4 , buf_splitterG5ton39n237_splitterG5ton236n237_1 , 0 , splitterG5ton236n237 );
splitter_AQFP splitterG6ton36n240_( clk_3 , G6 , 0 , splitterG6ton36n240 );
splitter_AQFP splitterG6ton156n240_( clk_5 , splitterG6ton36n240 , 0 , splitterG6ton156n240 );
splitter_AQFP splitterG6ton239n240_( clk_5 , buf_splitterG6ton156n240_splitterG6ton239n240_1 , 0 , splitterG6ton239n240 );
splitter_AQFP splitterG7ton36n243_( clk_3 , G7 , 0 , splitterG7ton36n243 );
splitter_AQFP splitterG7ton117n243_( clk_5 , splitterG7ton36n243 , 0 , splitterG7ton117n243 );
splitter_AQFP splitterG7ton242n243_( clk_5 , buf_splitterG7ton117n243_splitterG7ton242n243_1 , 0 , splitterG7ton242n243 );
splitter_AQFP splitterG8ton143n246_( clk_3 , G8 , 0 , splitterG8ton143n246 );
splitter_AQFP splitterG8ton144n246_( clk_5 , splitterG8ton143n246 , 0 , splitterG8ton144n246 );
splitter_AQFP splitterG8ton159n246_( clk_7 , splitterG8ton144n246 , 0 , splitterG8ton159n246 );
splitter_AQFP splitterG8ton245n246_( clk_5 , buf_splitterG8ton159n246_splitterG8ton245n246_1 , 0 , splitterG8ton245n246 );
splitter_AQFP splitterG9ton103n250_( clk_3 , G9 , 0 , splitterG9ton103n250 );
splitter_AQFP splitterG9ton58n250_( clk_7 , buf_splitterG9ton103n250_splitterG9ton58n250_1 , 0 , splitterG9ton58n250 );
splitter_AQFP splitterG9ton249n250_( clk_4 , buf_splitterG9ton58n250_splitterG9ton249n250_1 , 0 , splitterG9ton249n250 );
splitter_AQFP splitterfromn34_( clk_7 , n34 , 0 , splitterfromn34 );
splitter_AQFP splittern35ton269n252_( clk_4 , buf_n35_splittern35ton269n252_1 , 0 , splittern35ton269n252 );
splitter_AQFP splittern35ton78n252_( clk_6 , splittern35ton269n252 , 0 , splittern35ton78n252 );
splitter_AQFP splitterfromn38_( clk_6 , n38 , 0 , splitterfromn38 );
splitter_AQFP splittern41ton93n55_( clk_2 , n41 , 0 , splittern41ton93n55 );
splitter_AQFP splittern41ton54n55_( clk_3 , splittern41ton93n55 , 0 , splittern41ton54n55 );
splitter_AQFP splitterfromn44_( clk_1 , n44 , 0 , splitterfromn44 );
splitter_AQFP splitterfromn47_( clk_6 , n47 , 0 , splitterfromn47 );
splitter_AQFP splittern50ton51n187_( clk_1 , n50 , 0 , splittern50ton51n187 );
splitter_AQFP splitterfromn53_( clk_4 , n53 , 0 , splitterfromn53 );
splitter_AQFP splittern56ton70n299_( clk_7 , n56 , 0 , splittern56ton70n299 );
splitter_AQFP splitterfromn57_( clk_7 , n57 , 0 , splitterfromn57 );
splitter_AQFP splitterfromn60_( clk_2 , n60 , 0 , splitterfromn60 );
splitter_AQFP splittern63ton163n65_( clk_6 , n63 , 0 , splittern63ton163n65 );
splitter_AQFP splittern66ton85n68_( clk_1 , n66 , 0 , splittern66ton85n68 );
splitter_AQFP splitterfromn69_( clk_6 , n69 , 0 , splitterfromn69 );
splitter_AQFP splitterfromn72_( clk_2 , n72 , 0 , splitterfromn72 );
splitter_AQFP splittern73ton75n278_( clk_4 , n73 , 0 , splittern73ton75n278 );
splitter_AQFP splittern74ton75n275_( clk_3 , buf_n74_splittern74ton75n275_1 , 0 , splittern74ton75n275 );
splitter_AQFP splittern77ton271n253_( clk_7 , n77 , 0 , splittern77ton271n253 );
splitter_AQFP splitterfromn78_( clk_1 , n78 , 0 , splitterfromn78 );
splitter_AQFP splitterfromn81_( clk_6 , n81 , 0 , splitterfromn81 );
splitter_AQFP splitterfromn84_( clk_1 , n84 , 0 , splitterfromn84 );
splitter_AQFP splittern87ton189n97_( clk_4 , n87 , 0 , splittern87ton189n97 );
splitter_AQFP splittern87ton308n97_( clk_5 , splittern87ton189n97 , 0 , splittern87ton308n97 );
splitter_AQFP splitterfromn88_( clk_5 , n88 , 0 , splitterfromn88 );
splitter_AQFP splitterfromn89_( clk_7 , n89 , 0 , splitterfromn89 );
splitter_AQFP splitterfromn92_( clk_2 , n92 , 0 , splitterfromn92 );
splitter_AQFP splitterfromn95_( clk_5 , n95 , 0 , splitterfromn95 );
splitter_AQFP splitterfromn98_( clk_8 , n98 , 0 , splitterfromn98 );
splitter_AQFP splitterfromn99_( clk_2 , n99 , 0 , splitterfromn99 );
splitter_AQFP splittern105ton106n309_( clk_7 , n105 , 0 , splittern105ton106n309 );
splitter_AQFP splittern105ton308n309_( clk_4 , buf_splittern105ton106n309_splittern105ton308n309_1 , 0 , splittern105ton308n309 );
splitter_AQFP splittern108ton114n141_( clk_2 , n108 , 0 , splittern108ton114n141 );
splitter_AQFP splitterfromn109_( clk_5 , n109 , 0 , splitterfromn109 );
splitter_AQFP splitterfromn110_( clk_7 , n110 , 0 , splitterfromn110 );
splitter_AQFP splitterfromn113_( clk_2 , n113 , 0 , splitterfromn113 );
splitter_AQFP splitterfromn116_( clk_5 , n116 , 0 , splitterfromn116 );
splitter_AQFP splitterfromn119_( clk_1 , n119 , 0 , splitterfromn119 );
splitter_AQFP splitterfromn122_( clk_4 , n122 , 0 , splitterfromn122 );
splitter_AQFP splitterfromn125_( clk_8 , n125 , 0 , splitterfromn125 );
splitter_AQFP splitterfromn126_( clk_2 , n126 , 0 , splitterfromn126 );
splitter_AQFP splitterfromn127_( clk_7 , n127 , 0 , splitterfromn127 );
splitter_AQFP splittern128ton129n295_( clk_1 , buf_n128_splittern128ton129n295_1 , 0 , splittern128ton129n295 );
splitter_AQFP splitterfromn133_( clk_7 , n133 , 0 , splitterfromn133 );
splitter_AQFP splitterfromn136_( clk_6 , n136 , 0 , splitterfromn136 );
splitter_AQFP splitterfromn139_( clk_2 , n139 , 0 , splitterfromn139 );
splitter_AQFP splitterfromn142_( clk_5 , n142 , 0 , splitterfromn142 );
splitter_AQFP splitterfromn145_( clk_8 , n145 , 0 , splitterfromn145 );
splitter_AQFP splitterfromn148_( clk_4 , n148 , 0 , splitterfromn148 );
splitter_AQFP splitterfromn151_( clk_8 , n151 , 0 , splitterfromn151 );
splitter_AQFP splitterfromn152_( clk_2 , n152 , 0 , splitterfromn152 );
splitter_AQFP splitterfromn158_( clk_8 , n158 , 0 , splitterfromn158 );
splitter_AQFP splitterfromn161_( clk_3 , n161 , 0 , splitterfromn161 );
splitter_AQFP splitterfromn162_( clk_8 , n162 , 0 , splitterfromn162 );
splitter_AQFP splitterfromn165_( clk_1 , n165 , 0 , splitterfromn165 );
splitter_AQFP splitterfromn168_( clk_4 , n168 , 0 , splitterfromn168 );
splitter_AQFP splitterfromn171_( clk_8 , n171 , 0 , splitterfromn171 );
splitter_AQFP splitterfromn172_( clk_2 , n172 , 0 , splitterfromn172 );
splitter_AQFP splittern177ton197n272_( clk_7 , n177 , 0 , splittern177ton197n272 );
splitter_AQFP splittern178ton269n232_( clk_3 , buf_n178_splittern178ton269n232_1 , 0 , splittern178ton269n232 );
splitter_AQFP splittern178ton196n232_( clk_5 , splittern178ton269n232 , 0 , splittern178ton196n232 );
splitter_AQFP splitterfromn179_( clk_7 , n179 , 0 , splitterfromn179 );
splitter_AQFP splitterfromn182_( clk_7 , n182 , 0 , splitterfromn182 );
splitter_AQFP splitterfromn185_( clk_2 , n185 , 0 , splitterfromn185 );
splitter_AQFP splitterfromn188_( clk_5 , n188 , 0 , splitterfromn188 );
splitter_AQFP splitterfromn191_( clk_1 , n191 , 0 , splitterfromn191 );
splitter_AQFP splittern192ton193n284_( clk_3 , n192 , 0 , splittern192ton193n284 );
splitter_AQFP splittern195ton196n270_( clk_6 , n195 , 0 , splittern195ton196n270 );
splitter_AQFP splitterfromn197_( clk_1 , n197 , 0 , splitterfromn197 );
splitter_AQFP splitterfromn198_( clk_3 , n198 , 0 , splitterfromn198 );
splitter_AQFP splitterfromn199_( clk_7 , buf_n199_splitterfromn199_1 , 0 , splitterfromn199 );
splitter_AQFP splitterfromn200_( clk_1 , buf_n200_splitterfromn200_1 , 0 , splitterfromn200 );
splitter_AQFP splitterfromn201_( clk_4 , n201 , 0 , splitterfromn201 );
splitter_AQFP splittern203ton204n298_( clk_2 , n203 , 0 , splittern203ton204n298 );
splitter_AQFP splittern203ton321n298_( clk_5 , buf_splittern203ton204n298_splittern203ton321n298_1 , 0 , splittern203ton321n298 );
splitter_AQFP splittern203ton279n298_( clk_7 , splittern203ton321n298 , 0 , splittern203ton279n298 );
splitter_AQFP splittern203ton285n298_( clk_1 , splittern203ton279n298 , 0 , splittern203ton285n298 );
splitter_AQFP splitterfromn204_( clk_5 , n204 , 0 , splitterfromn204 );
splitter_AQFP splitterfromn205_( clk_2 , buf_n205_splitterfromn205_1 , 0 , splitterfromn205 );
splitter_AQFP splittern206ton267n217_( clk_5 , n206 , 0 , splittern206ton267n217 );
splitter_AQFP splittern206ton207n217_( clk_6 , splittern206ton267n217 , 0 , splittern206ton207n217 );
splitter_AQFP splittern206ton207n211_( clk_7 , splittern206ton207n217 , 0 , splittern206ton207n211 );
splitter_AQFP splittern206ton213n217_( clk_7 , splittern206ton207n217 , 0 , splittern206ton213n217 );
splitter_AQFP splitterfromn219_( clk_6 , buf_n219_splitterfromn219_1 , 0 , splitterfromn219 );
splitter_AQFP splittern221ton222n254_( clk_2 , buf_n221_splittern221ton222n254_1 , 0 , splittern221ton222n254 );
splitter_AQFP splittern222ton267n230_( clk_5 , n222 , 0 , splittern222ton267n230 );
splitter_AQFP splittern222ton223n230_( clk_6 , splittern222ton267n230 , 0 , splittern222ton223n230 );
splitter_AQFP splittern222ton226n230_( clk_7 , splittern222ton223n230 , 0 , splittern222ton226n230 );
splitter_AQFP splitterfromn234_( clk_3 , n234 , 0 , splitterfromn234 );
splitter_AQFP splittern235ton236n246_( clk_5 , n235 , 0 , splittern235ton236n246 );
splitter_AQFP splittern235ton239n240_( clk_6 , splittern235ton236n246 , 0 , splittern235ton239n240 );
splitter_AQFP splittern235ton242n246_( clk_6 , splittern235ton236n246 , 0 , splittern235ton242n246 );
splitter_AQFP splitterfromn248_( clk_5 , n248 , 0 , splitterfromn248 );
splitter_AQFP splittern254ton255n265_( clk_5 , n254 , 0 , splittern254ton255n265 );
splitter_AQFP splittern254ton255n259_( clk_6 , splittern254ton255n265 , 0 , splittern254ton255n259 );
splitter_AQFP splittern254ton261n265_( clk_6 , splittern254ton255n265 , 0 , splittern254ton261n265 );
splitter_AQFP splittern267ton275n320_( clk_7 , n267 , 0 , splittern267ton275n320 );
splitter_AQFP splittern267ton268n320_( clk_8 , splittern267ton275n320 , 0 , splittern267ton268n320 );
splitter_AQFP splitterfromn275_( clk_1 , n275 , 0 , splitterfromn275 );
splitter_AQFP splitterfromn281_( clk_1 , n281 , 0 , splitterfromn281 );
splitter_AQFP splitterfromn299_( clk_8 , buf_n299_splitterfromn299_1 , 0 , splitterfromn299 );
splitter_AQFP splitterfromn300_( clk_4 , buf_n300_splitterfromn300_1 , 0 , splitterfromn300 );
splitter_AQFP splitterfromn304_( clk_1 , n304 , 0 , splitterfromn304 );
splitter_AQFP splitterfromn311_( clk_8 , buf_n311_splitterfromn311_1 , 0 , splitterfromn311 );
splitter_AQFP splitterfromn312_( clk_4 , buf_n312_splitterfromn312_1 , 0 , splitterfromn312 );
splitter_AQFP splitterfromn316_( clk_1 , n316 , 0 , splitterfromn316 );

endmodule